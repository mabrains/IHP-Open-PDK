.SUBCKT LVL_LVMOS
MN1 D1 G1 S1 B sg13_hv_nmos w=0.6u l=0.45u ng=1 m=1 
MN2 D2 G2 S2 B sg13_hv_nmos w=0.8u l=0.45u ng=1 m=1 
MN3 D3 G3 S3 B sg13_hv_nmos w=0.8u l=0.5u  ng=1 m=1 
MN4 D4 G4 S4 B sg13_hv_nmos w=1.0u l=1.0u  ng=2 m=1 
.ENDS
