# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 13:19:48 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_256x16_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_256x16_c2_bm_bist 0 0 ;
  SIZE 419.95 BY 136.97 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.05 0 284.31 0.26 ;
    END
  END A_DIN[8]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.64 0 135.9 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.56 0 284.82 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.13 0 135.39 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 292.72 0 292.98 0.26 ;
    END
  END A_BM[8]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.97 0 127.23 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 291.345 0 291.605 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 128.345 0 128.605 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.91 0 277.17 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.78 0 143.04 0.26 ;
    END
  END A_DOUT[7]
  PIN B_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 286.6 0 286.86 0.26 ;
    END
  END B_DIN[8]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.09 0 133.35 0.26 ;
    END
  END B_DIN[7]
  PIN B_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 285.07 0 285.33 0.26 ;
    END
  END B_BIST_DIN[8]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.62 0 134.88 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 278.085 0 278.345 0.26 ;
    END
  END B_BM[8]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 141.605 0 141.865 0.26 ;
    END
  END B_BM[7]
  PIN B_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 279.615 0 279.875 0.26 ;
    END
  END B_BIST_BM[8]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 140.075 0 140.335 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.74 0 294 0.26 ;
    END
  END B_DOUT[8]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.95 0 126.21 0.26 ;
    END
  END B_DOUT[7]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 400.545 0 404.965 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 382.865 0 387.285 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.185 0 369.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.505 0 351.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.825 0 334.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 312.145 0 316.565 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.465 0 298.885 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 276.785 0 281.205 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 247.195 0 250.005 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 236.895 0 239.705 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 221.445 0 224.255 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 211.145 0 213.955 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 205.995 0 208.805 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.695 0 198.505 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 180.245 0 183.055 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.945 0 172.755 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.745 0 143.165 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.065 0 125.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.385 0 107.805 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.705 0 90.125 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 136.97 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.385 0 413.805 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 391.705 0 396.125 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.025 0 378.445 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 356.345 0 360.765 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 338.665 0 343.085 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 320.985 0 325.405 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 303.305 0 307.725 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.625 0 290.045 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 242.045 0 244.855 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 231.745 0 234.555 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 226.595 0 229.405 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.295 0 219.105 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.845 0 203.655 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.545 0 193.355 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 185.395 0 188.205 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.095 0 177.905 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 0 134.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 0 116.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 0 98.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 0 81.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.385 53.41 413.805 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 391.705 53.41 396.125 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.025 53.41 378.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 356.345 53.41 360.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 338.665 53.41 343.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 320.985 53.41 325.405 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 303.305 53.41 307.725 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.625 53.41 290.045 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 53.41 134.325 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 53.41 116.645 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 53.41 98.965 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 53.41 81.285 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 136.97 ;
    END
  END VDDARRAY!
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 301.73 0 301.99 0.26 ;
    END
  END A_DIN[9]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.96 0 118.22 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 302.24 0 302.5 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.45 0 117.71 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 310.4 0 310.66 0.26 ;
    END
  END A_BM[9]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.29 0 109.55 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 309.025 0 309.285 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.665 0 110.925 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.59 0 294.85 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.1 0 125.36 0.26 ;
    END
  END A_DOUT[6]
  PIN B_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.28 0 304.54 0.26 ;
    END
  END B_DIN[9]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.41 0 115.67 0.26 ;
    END
  END B_DIN[6]
  PIN B_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 302.75 0 303.01 0.26 ;
    END
  END B_BIST_DIN[9]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.94 0 117.2 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 295.765 0 296.025 0.26 ;
    END
  END B_BM[9]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.925 0 124.185 0.26 ;
    END
  END B_BM[6]
  PIN B_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 297.295 0 297.555 0.26 ;
    END
  END B_BIST_BM[9]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.395 0 122.655 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.42 0 311.68 0.26 ;
    END
  END B_DOUT[9]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.27 0 108.53 0.26 ;
    END
  END B_DOUT[6]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 319.41 0 319.67 0.26 ;
    END
  END A_DIN[10]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.28 0 100.54 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 319.92 0 320.18 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.77 0 100.03 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 328.08 0 328.34 0.26 ;
    END
  END A_BM[10]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 91.61 0 91.87 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 326.705 0 326.965 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 92.985 0 93.245 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 312.27 0 312.53 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 107.42 0 107.68 0.26 ;
    END
  END A_DOUT[5]
  PIN B_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 321.96 0 322.22 0.26 ;
    END
  END B_DIN[10]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 97.73 0 97.99 0.26 ;
    END
  END B_DIN[5]
  PIN B_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 320.43 0 320.69 0.26 ;
    END
  END B_BIST_DIN[10]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.26 0 99.52 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 313.445 0 313.705 0.26 ;
    END
  END B_BM[10]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 106.245 0 106.505 0.26 ;
    END
  END B_BM[5]
  PIN B_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 314.975 0 315.235 0.26 ;
    END
  END B_BIST_BM[10]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.715 0 104.975 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 329.1 0 329.36 0.26 ;
    END
  END B_DOUT[10]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 90.59 0 90.85 0.26 ;
    END
  END B_DOUT[5]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.09 0 337.35 0.26 ;
    END
  END A_DIN[11]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.6 0 82.86 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.6 0 337.86 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.09 0 82.35 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 345.76 0 346.02 0.26 ;
    END
  END A_BM[11]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 73.93 0 74.19 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 344.385 0 344.645 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 75.305 0 75.565 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 329.95 0 330.21 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.74 0 90 0.26 ;
    END
  END A_DOUT[4]
  PIN B_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.64 0 339.9 0.26 ;
    END
  END B_DIN[11]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 80.05 0 80.31 0.26 ;
    END
  END B_DIN[4]
  PIN B_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.11 0 338.37 0.26 ;
    END
  END B_BIST_DIN[11]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.58 0 81.84 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 331.125 0 331.385 0.26 ;
    END
  END B_BM[11]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.565 0 88.825 0.26 ;
    END
  END B_BM[4]
  PIN B_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 332.655 0 332.915 0.26 ;
    END
  END B_BIST_BM[11]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 87.035 0 87.295 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.78 0 347.04 0.26 ;
    END
  END B_DOUT[11]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.91 0 73.17 0.26 ;
    END
  END B_DOUT[4]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 354.77 0 355.03 0.26 ;
    END
  END A_DIN[12]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.28 0 355.54 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 363.44 0 363.7 0.26 ;
    END
  END A_BM[12]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.065 0 362.325 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.63 0 347.89 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 357.32 0 357.58 0.26 ;
    END
  END B_DIN[12]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.79 0 356.05 0.26 ;
    END
  END B_BIST_DIN[12]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 348.805 0 349.065 0.26 ;
    END
  END B_BM[12]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 350.335 0 350.595 0.26 ;
    END
  END B_BIST_BM[12]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.46 0 364.72 0.26 ;
    END
  END B_DOUT[12]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.45 0 372.71 0.26 ;
    END
  END A_DIN[13]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.96 0 373.22 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 381.12 0 381.38 0.26 ;
    END
  END A_BM[13]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.745 0 380.005 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 365.31 0 365.57 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 375 0 375.26 0.26 ;
    END
  END B_DIN[13]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.47 0 373.73 0.26 ;
    END
  END B_BIST_DIN[13]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 366.485 0 366.745 0.26 ;
    END
  END B_BM[13]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.015 0 368.275 0.26 ;
    END
  END B_BIST_BM[13]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.14 0 382.4 0.26 ;
    END
  END B_DOUT[13]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.13 0 390.39 0.26 ;
    END
  END A_DIN[14]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.64 0 390.9 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 398.8 0 399.06 0.26 ;
    END
  END A_BM[14]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 397.425 0 397.685 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.99 0 383.25 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 392.68 0 392.94 0.26 ;
    END
  END B_DIN[14]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 391.15 0 391.41 0.26 ;
    END
  END B_BIST_DIN[14]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.165 0 384.425 0.26 ;
    END
  END B_BM[14]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 385.695 0 385.955 0.26 ;
    END
  END B_BIST_BM[14]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 399.82 0 400.08 0.26 ;
    END
  END B_DOUT[14]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 407.81 0 408.07 0.26 ;
    END
  END A_DIN[15]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 408.32 0 408.58 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 416.48 0 416.74 0.26 ;
    END
  END A_BM[15]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 415.105 0 415.365 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.67 0 400.93 0.26 ;
    END
  END A_DOUT[15]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 410.36 0 410.62 0.26 ;
    END
  END B_DIN[15]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 408.83 0 409.09 0.26 ;
    END
  END B_BIST_DIN[15]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.845 0 402.105 0.26 ;
    END
  END B_BM[15]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 403.375 0 403.635 0.26 ;
    END
  END B_BIST_BM[15]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 417.5 0 417.76 0.26 ;
    END
  END B_DOUT[15]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.065 0 226.325 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.675 0 231.935 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.625 0 193.885 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.015 0 188.275 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.575 0 226.835 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.185 0 232.445 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.115 0 193.375 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 187.505 0 187.765 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 235.245 0 235.505 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 235.755 0 236.015 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 184.445 0 184.705 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 183.935 0 184.195 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 234.225 0 234.485 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 234.735 0 234.995 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 185.465 0 185.725 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 184.955 0 185.215 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.845 0 215.105 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.355 0 215.615 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.845 0 205.105 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.335 0 204.595 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.825 0 214.085 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.335 0 214.595 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.865 0 206.125 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.355 0 205.615 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 237.795 0 238.055 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 237.285 0 237.545 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.895 0 182.155 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.405 0 182.665 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 236.775 0 237.035 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 236.265 0 236.525 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.915 0 183.175 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 183.425 0 183.685 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.535 0 224.795 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.105 0 228.365 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.595 0 227.855 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 225.045 0 225.305 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 245.445 0 245.705 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.155 0 195.415 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 191.585 0 191.845 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.095 0 192.355 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 194.645 0 194.905 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 174.245 0 174.505 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 150.4115 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 15.73 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.733454 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.085 0 227.345 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.005 0 223.265 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 229.635 0 229.895 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 229.125 0 229.385 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.515 0 223.775 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 150.9886 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 15.73 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.770142 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.605 0 192.865 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.685 0 196.945 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 190.055 0 190.315 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 190.565 0 190.825 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.175 0 196.435 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 419.95 136.97 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 136.94 ;
      RECT 1.135 136.21 1.335 136.94 ;
      RECT 1.545 136.21 1.905 136.94 ;
      RECT 2.115 136.21 2.315 136.94 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 136.21 2.97 136.94 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 136.21 3.54 136.94 ;
      RECT 3.835 136.21 4.035 136.94 ;
      RECT 4.33 136.21 4.69 136.94 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 136.21 5.1 136.94 ;
      RECT 5.555 136.21 5.755 136.94 ;
      RECT 5.965 136.21 6.325 136.94 ;
      RECT 6.535 136.21 6.735 136.94 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 136.21 7.39 136.94 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 136.21 7.96 136.94 ;
      RECT 8.255 136.21 8.455 136.94 ;
      RECT 8.75 136.21 9.11 136.94 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 136.21 9.52 136.94 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 136.21 10.175 136.94 ;
      RECT 10.385 136.21 10.745 136.94 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 136.21 11.155 136.94 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 136.21 11.81 136.94 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 136.21 12.38 136.94 ;
      RECT 12.675 136.21 12.875 136.94 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 136.21 13.53 136.94 ;
      RECT 13.74 136.21 13.94 136.94 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 136.21 14.595 136.94 ;
      RECT 14.805 136.21 15.165 136.94 ;
      RECT 15.375 136.21 15.575 136.94 ;
      RECT 16.03 136.21 16.23 136.94 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 136.21 16.8 136.94 ;
      RECT 17.095 136.21 17.295 136.94 ;
      RECT 17.59 136.21 17.95 136.94 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 136.21 18.36 136.94 ;
      RECT 18.815 136.21 19.015 136.94 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 136.21 19.585 136.94 ;
      RECT 19.795 136.21 19.995 136.94 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 136.21 20.65 136.94 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 136.21 21.22 136.94 ;
      RECT 21.515 136.21 21.715 136.94 ;
      RECT 22.01 136.21 22.37 136.94 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 136.21 22.78 136.94 ;
      RECT 23.235 136.21 23.435 136.94 ;
      RECT 23.645 136.21 24.005 136.94 ;
      RECT 24.215 136.21 24.415 136.94 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 136.21 25.07 136.94 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 136.21 25.64 136.94 ;
      RECT 25.935 136.21 26.135 136.94 ;
      RECT 26.43 136.21 26.79 136.94 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 136.21 27.2 136.94 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 136.21 27.855 136.94 ;
      RECT 28.065 136.21 28.425 136.94 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 136.21 28.835 136.94 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 136.21 29.49 136.94 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 136.21 30.06 136.94 ;
      RECT 30.355 136.21 30.555 136.94 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 136.21 31.21 136.94 ;
      RECT 31.42 136.21 31.62 136.94 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 136.21 32.275 136.94 ;
      RECT 32.485 136.21 32.845 136.94 ;
      RECT 33.055 136.21 33.255 136.94 ;
      RECT 33.71 136.21 33.91 136.94 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 136.21 34.48 136.94 ;
      RECT 34.775 136.21 34.975 136.94 ;
      RECT 35.27 136.21 35.63 136.94 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 136.21 36.04 136.94 ;
      RECT 36.495 136.21 36.695 136.94 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 136.21 37.265 136.94 ;
      RECT 37.475 136.21 37.675 136.94 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 136.21 38.33 136.94 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 136.21 38.9 136.94 ;
      RECT 39.195 136.21 39.395 136.94 ;
      RECT 39.69 136.21 40.05 136.94 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 136.21 40.46 136.94 ;
      RECT 40.915 136.21 41.115 136.94 ;
      RECT 41.325 136.21 41.685 136.94 ;
      RECT 41.895 136.21 42.095 136.94 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 136.21 42.75 136.94 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 136.21 43.32 136.94 ;
      RECT 43.615 136.21 43.815 136.94 ;
      RECT 44.11 136.21 44.47 136.94 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 136.21 44.88 136.94 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 136.21 45.535 136.94 ;
      RECT 45.745 136.21 46.105 136.94 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 136.21 46.515 136.94 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 136.21 47.17 136.94 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 136.21 47.74 136.94 ;
      RECT 48.035 136.21 48.235 136.94 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 136.21 48.89 136.94 ;
      RECT 49.1 136.21 49.3 136.94 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 136.21 49.955 136.94 ;
      RECT 50.165 136.21 50.525 136.94 ;
      RECT 50.735 136.21 50.935 136.94 ;
      RECT 51.39 136.21 51.59 136.94 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 136.21 52.16 136.94 ;
      RECT 52.455 136.21 52.655 136.94 ;
      RECT 52.95 136.21 53.31 136.94 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 136.21 53.72 136.94 ;
      RECT 54.175 136.21 54.375 136.94 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 136.21 54.945 136.94 ;
      RECT 55.155 136.21 55.355 136.94 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 136.21 56.01 136.94 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 136.21 56.58 136.94 ;
      RECT 56.875 136.21 57.075 136.94 ;
      RECT 57.37 136.21 57.73 136.94 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 136.21 58.14 136.94 ;
      RECT 58.595 136.21 58.795 136.94 ;
      RECT 59.005 136.21 59.365 136.94 ;
      RECT 59.575 136.21 59.775 136.94 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 136.21 60.43 136.94 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 136.21 61 136.94 ;
      RECT 61.295 136.21 61.495 136.94 ;
      RECT 61.79 136.21 62.15 136.94 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 136.21 62.56 136.94 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 136.21 63.215 136.94 ;
      RECT 63.425 136.21 63.785 136.94 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 136.21 64.195 136.94 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 136.21 64.85 136.94 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 136.21 65.42 136.94 ;
      RECT 65.715 136.21 65.915 136.94 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 136.21 66.57 136.94 ;
      RECT 66.78 136.21 66.98 136.94 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 136.21 67.635 136.94 ;
      RECT 67.845 136.21 68.205 136.94 ;
      RECT 68.415 136.21 68.615 136.94 ;
      RECT 69.07 136.21 69.27 136.94 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 136.21 69.84 136.94 ;
      RECT 70.135 136.21 70.335 136.94 ;
      RECT 70.63 136.21 70.99 136.94 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 136.21 71.4 136.94 ;
      RECT 71.855 136.21 72.055 136.94 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 72.265 136.21 72.625 136.94 ;
      RECT 72.835 136.21 73.035 136.94 ;
      RECT 72.91 0.52 73.17 7.78 ;
      RECT 73.42 0.3 73.68 5.235 ;
      RECT 73.49 136.21 73.69 136.94 ;
      RECT 73.93 0.52 74.19 5.57 ;
      RECT 73.9 136.21 74.26 136.94 ;
      RECT 74.555 136.21 74.755 136.94 ;
      RECT 75.05 136.21 75.41 136.94 ;
      RECT 75.305 0.52 75.565 6.28 ;
      RECT 75.62 136.21 75.82 136.94 ;
      RECT 76.275 136.21 76.475 136.94 ;
      RECT 76.685 136.21 77.045 136.94 ;
      RECT 77.255 136.21 77.455 136.94 ;
      RECT 76.99 0.18 77.76 0.88 ;
      RECT 77.91 136.21 78.11 136.94 ;
      RECT 78.01 0.3 78.27 8.7 ;
      RECT 78.32 136.21 78.68 136.94 ;
      RECT 78.975 136.21 79.175 136.94 ;
      RECT 79.47 136.21 79.83 136.94 ;
      RECT 80.56 0.155 81.33 0.445 ;
      RECT 80.56 0.155 80.82 8.665 ;
      RECT 81.07 0.155 81.33 8.665 ;
      RECT 80.04 136.21 80.24 136.94 ;
      RECT 80.05 0.52 80.31 9.955 ;
      RECT 80.695 136.21 80.895 136.94 ;
      RECT 81.105 136.21 81.465 136.94 ;
      RECT 81.58 0.52 81.84 11.315 ;
      RECT 81.675 136.21 81.875 136.94 ;
      RECT 82.09 0.52 82.35 13.45 ;
      RECT 82.33 136.21 82.53 136.94 ;
      RECT 82.6 0.52 82.86 14.115 ;
      RECT 82.74 136.21 83.1 136.94 ;
      RECT 83.395 136.21 83.595 136.94 ;
      RECT 84.795 0.155 85.565 0.445 ;
      RECT 84.795 0.155 85.055 13.21 ;
      RECT 85.305 0.155 85.565 13.21 ;
      RECT 83.89 136.21 84.25 136.94 ;
      RECT 84.46 136.21 84.66 136.94 ;
      RECT 85.815 0.18 86.585 0.88 ;
      RECT 85.815 0.18 86.075 12.9 ;
      RECT 86.325 0.18 86.585 12.9 ;
      RECT 85.115 136.21 85.315 136.94 ;
      RECT 85.525 136.21 85.885 136.94 ;
      RECT 86.095 136.21 86.295 136.94 ;
      RECT 86.75 136.21 86.95 136.94 ;
      RECT 87.035 0.52 87.295 2.82 ;
      RECT 87.16 136.21 87.52 136.94 ;
      RECT 87.815 136.21 88.015 136.94 ;
      RECT 88.31 136.21 88.67 136.94 ;
      RECT 88.565 0.52 88.825 2.82 ;
      RECT 88.88 136.21 89.08 136.94 ;
      RECT 89.535 136.21 89.735 136.94 ;
      RECT 89.74 0.52 90 4.315 ;
      RECT 89.945 136.21 90.305 136.94 ;
      RECT 90.515 136.21 90.715 136.94 ;
      RECT 90.59 0.52 90.85 7.78 ;
      RECT 91.1 0.3 91.36 5.235 ;
      RECT 91.17 136.21 91.37 136.94 ;
      RECT 91.61 0.52 91.87 5.57 ;
      RECT 91.58 136.21 91.94 136.94 ;
      RECT 92.235 136.21 92.435 136.94 ;
      RECT 92.73 136.21 93.09 136.94 ;
      RECT 92.985 0.52 93.245 6.28 ;
      RECT 93.3 136.21 93.5 136.94 ;
      RECT 93.955 136.21 94.155 136.94 ;
      RECT 94.365 136.21 94.725 136.94 ;
      RECT 94.935 136.21 95.135 136.94 ;
      RECT 94.67 0.18 95.44 0.88 ;
      RECT 95.59 136.21 95.79 136.94 ;
      RECT 95.69 0.3 95.95 8.7 ;
      RECT 96 136.21 96.36 136.94 ;
      RECT 96.655 136.21 96.855 136.94 ;
      RECT 97.15 136.21 97.51 136.94 ;
      RECT 98.24 0.155 99.01 0.445 ;
      RECT 98.24 0.155 98.5 8.665 ;
      RECT 98.75 0.155 99.01 8.665 ;
      RECT 97.72 136.21 97.92 136.94 ;
      RECT 97.73 0.52 97.99 9.955 ;
      RECT 98.375 136.21 98.575 136.94 ;
      RECT 98.785 136.21 99.145 136.94 ;
      RECT 99.26 0.52 99.52 11.315 ;
      RECT 99.355 136.21 99.555 136.94 ;
      RECT 99.77 0.52 100.03 13.45 ;
      RECT 100.01 136.21 100.21 136.94 ;
      RECT 100.28 0.52 100.54 14.115 ;
      RECT 100.42 136.21 100.78 136.94 ;
      RECT 101.075 136.21 101.275 136.94 ;
      RECT 102.475 0.155 103.245 0.445 ;
      RECT 102.475 0.155 102.735 13.21 ;
      RECT 102.985 0.155 103.245 13.21 ;
      RECT 101.57 136.21 101.93 136.94 ;
      RECT 102.14 136.21 102.34 136.94 ;
      RECT 103.495 0.18 104.265 0.88 ;
      RECT 103.495 0.18 103.755 12.9 ;
      RECT 104.005 0.18 104.265 12.9 ;
      RECT 102.795 136.21 102.995 136.94 ;
      RECT 103.205 136.21 103.565 136.94 ;
      RECT 103.775 136.21 103.975 136.94 ;
      RECT 104.43 136.21 104.63 136.94 ;
      RECT 104.715 0.52 104.975 2.82 ;
      RECT 104.84 136.21 105.2 136.94 ;
      RECT 105.495 136.21 105.695 136.94 ;
      RECT 105.99 136.21 106.35 136.94 ;
      RECT 106.245 0.52 106.505 2.82 ;
      RECT 106.56 136.21 106.76 136.94 ;
      RECT 107.215 136.21 107.415 136.94 ;
      RECT 107.42 0.52 107.68 4.315 ;
      RECT 107.625 136.21 107.985 136.94 ;
      RECT 108.195 136.21 108.395 136.94 ;
      RECT 108.27 0.52 108.53 7.78 ;
      RECT 108.78 0.3 109.04 5.235 ;
      RECT 108.85 136.21 109.05 136.94 ;
      RECT 109.29 0.52 109.55 5.57 ;
      RECT 109.26 136.21 109.62 136.94 ;
      RECT 109.915 136.21 110.115 136.94 ;
      RECT 110.41 136.21 110.77 136.94 ;
      RECT 110.665 0.52 110.925 6.28 ;
      RECT 110.98 136.21 111.18 136.94 ;
      RECT 111.635 136.21 111.835 136.94 ;
      RECT 112.045 136.21 112.405 136.94 ;
      RECT 112.615 136.21 112.815 136.94 ;
      RECT 112.35 0.18 113.12 0.88 ;
      RECT 113.27 136.21 113.47 136.94 ;
      RECT 113.37 0.3 113.63 8.7 ;
      RECT 113.68 136.21 114.04 136.94 ;
      RECT 114.335 136.21 114.535 136.94 ;
      RECT 114.83 136.21 115.19 136.94 ;
      RECT 115.92 0.155 116.69 0.445 ;
      RECT 115.92 0.155 116.18 8.665 ;
      RECT 116.43 0.155 116.69 8.665 ;
      RECT 115.4 136.21 115.6 136.94 ;
      RECT 115.41 0.52 115.67 9.955 ;
      RECT 116.055 136.21 116.255 136.94 ;
      RECT 116.465 136.21 116.825 136.94 ;
      RECT 116.94 0.52 117.2 11.315 ;
      RECT 117.035 136.21 117.235 136.94 ;
      RECT 117.45 0.52 117.71 13.45 ;
      RECT 117.69 136.21 117.89 136.94 ;
      RECT 117.96 0.52 118.22 14.115 ;
      RECT 118.1 136.21 118.46 136.94 ;
      RECT 118.755 136.21 118.955 136.94 ;
      RECT 120.155 0.155 120.925 0.445 ;
      RECT 120.155 0.155 120.415 13.21 ;
      RECT 120.665 0.155 120.925 13.21 ;
      RECT 119.25 136.21 119.61 136.94 ;
      RECT 119.82 136.21 120.02 136.94 ;
      RECT 121.175 0.18 121.945 0.88 ;
      RECT 121.175 0.18 121.435 12.9 ;
      RECT 121.685 0.18 121.945 12.9 ;
      RECT 120.475 136.21 120.675 136.94 ;
      RECT 120.885 136.21 121.245 136.94 ;
      RECT 121.455 136.21 121.655 136.94 ;
      RECT 122.11 136.21 122.31 136.94 ;
      RECT 122.395 0.52 122.655 2.82 ;
      RECT 122.52 136.21 122.88 136.94 ;
      RECT 123.175 136.21 123.375 136.94 ;
      RECT 123.67 136.21 124.03 136.94 ;
      RECT 123.925 0.52 124.185 2.82 ;
      RECT 124.24 136.21 124.44 136.94 ;
      RECT 124.895 136.21 125.095 136.94 ;
      RECT 125.1 0.52 125.36 4.315 ;
      RECT 125.305 136.21 125.665 136.94 ;
      RECT 125.875 136.21 126.075 136.94 ;
      RECT 125.95 0.52 126.21 7.78 ;
      RECT 126.46 0.3 126.72 5.235 ;
      RECT 126.53 136.21 126.73 136.94 ;
      RECT 126.97 0.52 127.23 5.57 ;
      RECT 126.94 136.21 127.3 136.94 ;
      RECT 127.595 136.21 127.795 136.94 ;
      RECT 128.09 136.21 128.45 136.94 ;
      RECT 128.345 0.52 128.605 6.28 ;
      RECT 128.66 136.21 128.86 136.94 ;
      RECT 129.315 136.21 129.515 136.94 ;
      RECT 129.725 136.21 130.085 136.94 ;
      RECT 130.295 136.21 130.495 136.94 ;
      RECT 130.03 0.18 130.8 0.88 ;
      RECT 130.95 136.21 131.15 136.94 ;
      RECT 131.05 0.3 131.31 8.7 ;
      RECT 131.36 136.21 131.72 136.94 ;
      RECT 132.015 136.21 132.215 136.94 ;
      RECT 132.51 136.21 132.87 136.94 ;
      RECT 133.6 0.155 134.37 0.445 ;
      RECT 133.6 0.155 133.86 8.665 ;
      RECT 134.11 0.155 134.37 8.665 ;
      RECT 133.08 136.21 133.28 136.94 ;
      RECT 133.09 0.52 133.35 9.955 ;
      RECT 133.735 136.21 133.935 136.94 ;
      RECT 134.145 136.21 134.505 136.94 ;
      RECT 134.62 0.52 134.88 11.315 ;
      RECT 134.715 136.21 134.915 136.94 ;
      RECT 135.13 0.52 135.39 13.45 ;
      RECT 135.37 136.21 135.57 136.94 ;
      RECT 135.64 0.52 135.9 14.115 ;
      RECT 135.78 136.21 136.14 136.94 ;
      RECT 136.435 136.21 136.635 136.94 ;
      RECT 137.835 0.155 138.605 0.445 ;
      RECT 137.835 0.155 138.095 13.21 ;
      RECT 138.345 0.155 138.605 13.21 ;
      RECT 136.93 136.21 137.29 136.94 ;
      RECT 137.5 136.21 137.7 136.94 ;
      RECT 138.855 0.18 139.625 0.88 ;
      RECT 138.855 0.18 139.115 12.9 ;
      RECT 139.365 0.18 139.625 12.9 ;
      RECT 138.155 136.21 138.355 136.94 ;
      RECT 138.565 136.21 138.925 136.94 ;
      RECT 139.135 136.21 139.335 136.94 ;
      RECT 139.79 136.21 139.99 136.94 ;
      RECT 140.075 0.52 140.335 2.82 ;
      RECT 140.2 136.21 140.56 136.94 ;
      RECT 140.855 136.21 141.055 136.94 ;
      RECT 141.35 136.21 141.71 136.94 ;
      RECT 141.605 0.52 141.865 2.82 ;
      RECT 141.92 136.21 142.12 136.94 ;
      RECT 142.575 136.21 142.775 136.94 ;
      RECT 142.78 0.52 143.04 4.315 ;
      RECT 144.31 0.17 145.08 0.43 ;
      RECT 144.31 0.17 144.57 8.7 ;
      RECT 144.82 0.17 145.08 8.7 ;
      RECT 145.33 0.18 146.1 0.88 ;
      RECT 145.33 0.18 145.59 8.7 ;
      RECT 145.84 0.18 146.1 8.7 ;
      RECT 146.35 0.17 147.12 0.43 ;
      RECT 146.35 0.17 146.61 8.7 ;
      RECT 146.86 0.17 147.12 8.7 ;
      RECT 147.37 0.18 148.14 0.88 ;
      RECT 147.37 0.18 147.63 8.7 ;
      RECT 147.88 0.18 148.14 8.7 ;
      RECT 148.39 0.17 149.16 0.43 ;
      RECT 148.39 0.17 148.65 8.7 ;
      RECT 148.9 0.17 149.16 8.7 ;
      RECT 149.41 0.18 150.18 0.88 ;
      RECT 149.41 0.18 149.67 8.7 ;
      RECT 149.92 0.18 150.18 8.7 ;
      RECT 150.43 0.17 151.2 0.43 ;
      RECT 150.43 0.17 150.69 8.7 ;
      RECT 150.94 0.17 151.2 8.7 ;
      RECT 151.45 0.18 152.22 0.88 ;
      RECT 151.45 0.18 151.71 8.7 ;
      RECT 151.96 0.18 152.22 8.7 ;
      RECT 152.47 0.17 153.24 0.43 ;
      RECT 152.47 0.17 152.73 8.7 ;
      RECT 152.98 0.17 153.24 8.7 ;
      RECT 153.49 0.18 154.26 0.88 ;
      RECT 153.49 0.18 153.75 8.7 ;
      RECT 154 0.18 154.26 8.7 ;
      RECT 154.51 0.17 155.28 0.43 ;
      RECT 154.51 0.17 154.77 8.7 ;
      RECT 155.02 0.17 155.28 8.7 ;
      RECT 155.53 0.18 156.3 0.88 ;
      RECT 155.53 0.18 155.79 8.7 ;
      RECT 156.04 0.18 156.3 8.7 ;
      RECT 156.55 0.17 157.32 0.43 ;
      RECT 156.55 0.17 156.81 8.7 ;
      RECT 157.06 0.17 157.32 8.7 ;
      RECT 157.57 0.18 158.34 0.88 ;
      RECT 157.57 0.18 157.83 8.7 ;
      RECT 158.08 0.18 158.34 8.7 ;
      RECT 158.59 0.17 159.36 0.43 ;
      RECT 158.59 0.17 158.85 8.7 ;
      RECT 159.1 0.17 159.36 8.7 ;
      RECT 159.61 0.18 160.38 0.88 ;
      RECT 159.61 0.18 159.87 8.7 ;
      RECT 160.12 0.18 160.38 8.7 ;
      RECT 160.63 0.17 161.4 0.43 ;
      RECT 160.63 0.17 160.89 8.7 ;
      RECT 161.14 0.17 161.4 8.7 ;
      RECT 161.65 0.18 162.42 0.88 ;
      RECT 161.65 0.18 161.91 8.7 ;
      RECT 162.16 0.18 162.42 8.7 ;
      RECT 162.67 0.17 163.44 0.43 ;
      RECT 162.67 0.17 162.93 8.7 ;
      RECT 163.18 0.17 163.44 8.7 ;
      RECT 163.69 0.18 164.46 0.88 ;
      RECT 163.69 0.18 163.95 8.7 ;
      RECT 164.2 0.18 164.46 8.7 ;
      RECT 164.71 0.17 165.48 0.43 ;
      RECT 164.71 0.17 164.97 8.7 ;
      RECT 165.22 0.17 165.48 8.7 ;
      RECT 165.73 0.18 166.5 0.88 ;
      RECT 165.73 0.18 165.99 8.7 ;
      RECT 166.24 0.18 166.5 8.7 ;
      RECT 166.75 0.17 167.52 0.43 ;
      RECT 166.75 0.17 167.01 8.7 ;
      RECT 167.26 0.17 167.52 8.7 ;
      RECT 167.77 0.18 168.54 0.88 ;
      RECT 167.77 0.18 168.03 8.7 ;
      RECT 168.28 0.18 168.54 8.7 ;
      RECT 142.985 136.21 143.345 136.94 ;
      RECT 143.555 136.21 143.755 136.94 ;
      RECT 170.165 0.18 170.935 0.88 ;
      RECT 170.165 0.18 170.425 8.7 ;
      RECT 170.675 0.18 170.935 8.7 ;
      RECT 171.185 0.17 171.955 0.43 ;
      RECT 171.185 0.17 171.445 8.7 ;
      RECT 171.695 0.17 171.955 8.7 ;
      RECT 144.38 136.13 144.58 136.94 ;
      RECT 169.145 0.3 169.405 8.7 ;
      RECT 173.225 0.18 173.995 0.88 ;
      RECT 173.225 0.18 173.485 8.7 ;
      RECT 173.735 0.18 173.995 8.7 ;
      RECT 169.655 0.3 169.915 8.7 ;
      RECT 172.205 0 172.465 8.7 ;
      RECT 172.715 0 172.975 8.7 ;
      RECT 174.245 0.52 174.505 8.7 ;
      RECT 174.755 0.3 175.015 8.7 ;
      RECT 175.265 0.3 175.525 8.7 ;
      RECT 175.775 0.3 176.035 8.7 ;
      RECT 176.285 0.3 176.545 8.7 ;
      RECT 176.795 0.3 177.055 8.7 ;
      RECT 177.305 0.3 177.565 8.7 ;
      RECT 177.815 0.3 178.075 8.7 ;
      RECT 179.855 0.18 180.625 0.88 ;
      RECT 179.855 0.18 180.115 8.7 ;
      RECT 180.365 0.18 180.625 8.7 ;
      RECT 178.325 0.3 178.585 8.7 ;
      RECT 178.835 0 179.095 8.7 ;
      RECT 179.345 0 179.605 8.7 ;
      RECT 180.875 0 181.135 8.7 ;
      RECT 181.385 0 181.645 8.7 ;
      RECT 181.895 0.52 182.155 8.7 ;
      RECT 182.405 0.52 182.665 8.7 ;
      RECT 182.915 0.52 183.175 8.7 ;
      RECT 183.425 0.52 183.685 8.7 ;
      RECT 183.935 0.52 184.195 8.7 ;
      RECT 184.445 0.52 184.705 8.7 ;
      RECT 184.955 0.52 185.215 8.7 ;
      RECT 185.465 0.52 185.725 8.7 ;
      RECT 185.975 0.3 186.235 8.7 ;
      RECT 186.485 0.3 186.745 8.7 ;
      RECT 186.995 0.3 187.255 8.7 ;
      RECT 187.505 0.52 187.765 8.7 ;
      RECT 188.015 0.52 188.275 8.7 ;
      RECT 188.525 0.3 188.785 8.7 ;
      RECT 189.035 0.3 189.295 8.7 ;
      RECT 189.545 0.3 189.805 8.7 ;
      RECT 190.055 0.52 190.315 8.7 ;
      RECT 190.565 0.52 190.825 8.7 ;
      RECT 191.075 0.3 191.335 8.7 ;
      RECT 191.585 0.52 191.845 8.7 ;
      RECT 192.095 0.52 192.355 8.7 ;
      RECT 192.605 0.52 192.865 8.7 ;
      RECT 193.115 0.52 193.375 8.7 ;
      RECT 193.625 0.52 193.885 8.7 ;
      RECT 194.135 0.3 194.395 8.7 ;
      RECT 194.645 0.52 194.905 8.7 ;
      RECT 195.155 0.52 195.415 8.7 ;
      RECT 195.665 0.3 195.925 8.7 ;
      RECT 196.175 0.52 196.435 8.7 ;
      RECT 198.215 0.17 198.985 0.43 ;
      RECT 198.215 0.17 198.475 8.7 ;
      RECT 198.725 0.17 198.985 8.7 ;
      RECT 196.685 0.52 196.945 8.7 ;
      RECT 197.195 0.3 197.455 8.7 ;
      RECT 197.705 0.3 197.965 8.7 ;
      RECT 200.765 0.17 201.535 0.43 ;
      RECT 200.765 0.17 201.025 8.7 ;
      RECT 201.275 0.17 201.535 8.7 ;
      RECT 199.235 0.3 199.495 8.7 ;
      RECT 202.295 0.18 203.065 0.88 ;
      RECT 202.295 0.18 202.555 8.7 ;
      RECT 202.805 0.18 203.065 8.7 ;
      RECT 199.745 0.3 200.005 8.7 ;
      RECT 200.255 0.3 200.515 8.7 ;
      RECT 201.785 0.3 202.045 8.7 ;
      RECT 203.315 0 203.575 8.7 ;
      RECT 203.825 0 204.085 8.7 ;
      RECT 204.335 0.52 204.595 8.7 ;
      RECT 204.845 0.52 205.105 8.7 ;
      RECT 205.355 0.52 205.615 8.7 ;
      RECT 205.865 0.52 206.125 8.7 ;
      RECT 206.375 0 206.635 8.7 ;
      RECT 206.885 0 207.145 8.7 ;
      RECT 207.395 0.3 207.655 8.7 ;
      RECT 207.905 0.3 208.165 8.7 ;
      RECT 208.415 0 208.675 8.7 ;
      RECT 208.925 0 209.185 8.7 ;
      RECT 209.435 0.3 209.695 8.7 ;
      RECT 210.255 0.3 210.515 8.7 ;
      RECT 210.765 0 211.025 8.7 ;
      RECT 211.275 0 211.535 8.7 ;
      RECT 211.785 0.3 212.045 8.7 ;
      RECT 212.295 0.3 212.555 8.7 ;
      RECT 212.805 0 213.065 8.7 ;
      RECT 213.315 0 213.575 8.7 ;
      RECT 213.825 0.52 214.085 8.7 ;
      RECT 214.335 0.52 214.595 8.7 ;
      RECT 214.845 0.52 215.105 8.7 ;
      RECT 216.885 0.18 217.655 0.88 ;
      RECT 216.885 0.18 217.145 8.7 ;
      RECT 217.395 0.18 217.655 8.7 ;
      RECT 215.355 0.52 215.615 8.7 ;
      RECT 218.415 0.17 219.185 0.43 ;
      RECT 218.415 0.17 218.675 8.7 ;
      RECT 218.925 0.17 219.185 8.7 ;
      RECT 215.865 0 216.125 8.7 ;
      RECT 216.375 0 216.635 8.7 ;
      RECT 217.905 0.3 218.165 8.7 ;
      RECT 220.965 0.17 221.735 0.43 ;
      RECT 220.965 0.17 221.225 8.7 ;
      RECT 221.475 0.17 221.735 8.7 ;
      RECT 219.435 0.3 219.695 8.7 ;
      RECT 219.945 0.3 220.205 8.7 ;
      RECT 220.455 0.3 220.715 8.7 ;
      RECT 221.985 0.3 222.245 8.7 ;
      RECT 222.495 0.3 222.755 8.7 ;
      RECT 223.005 0.52 223.265 8.7 ;
      RECT 223.515 0.52 223.775 8.7 ;
      RECT 224.025 0.3 224.285 8.7 ;
      RECT 224.535 0.52 224.795 8.7 ;
      RECT 225.045 0.52 225.305 8.7 ;
      RECT 225.555 0.3 225.815 8.7 ;
      RECT 226.065 0.52 226.325 8.7 ;
      RECT 226.575 0.52 226.835 8.7 ;
      RECT 227.085 0.52 227.345 8.7 ;
      RECT 227.595 0.52 227.855 8.7 ;
      RECT 228.105 0.52 228.365 8.7 ;
      RECT 228.615 0.3 228.875 8.7 ;
      RECT 229.125 0.52 229.385 8.7 ;
      RECT 229.635 0.52 229.895 8.7 ;
      RECT 230.145 0.3 230.405 8.7 ;
      RECT 230.655 0.3 230.915 8.7 ;
      RECT 231.165 0.3 231.425 8.7 ;
      RECT 231.675 0.52 231.935 8.7 ;
      RECT 232.185 0.52 232.445 8.7 ;
      RECT 232.695 0.3 232.955 8.7 ;
      RECT 233.205 0.3 233.465 8.7 ;
      RECT 233.715 0.3 233.975 8.7 ;
      RECT 234.225 0.52 234.485 8.7 ;
      RECT 234.735 0.52 234.995 8.7 ;
      RECT 235.245 0.52 235.505 8.7 ;
      RECT 235.755 0.52 236.015 8.7 ;
      RECT 236.265 0.52 236.525 8.7 ;
      RECT 236.775 0.52 237.035 8.7 ;
      RECT 237.285 0.52 237.545 8.7 ;
      RECT 239.325 0.18 240.095 0.88 ;
      RECT 239.325 0.18 239.585 8.7 ;
      RECT 239.835 0.18 240.095 8.7 ;
      RECT 237.795 0.52 238.055 8.7 ;
      RECT 238.305 0 238.565 8.7 ;
      RECT 238.815 0 239.075 8.7 ;
      RECT 240.345 0 240.605 8.7 ;
      RECT 240.855 0 241.115 8.7 ;
      RECT 241.365 0.3 241.625 8.7 ;
      RECT 241.875 0.3 242.135 8.7 ;
      RECT 242.385 0.3 242.645 8.7 ;
      RECT 242.895 0.3 243.155 8.7 ;
      RECT 243.405 0.3 243.665 8.7 ;
      RECT 243.915 0.3 244.175 8.7 ;
      RECT 245.955 0.18 246.725 0.88 ;
      RECT 245.955 0.18 246.215 8.7 ;
      RECT 246.465 0.18 246.725 8.7 ;
      RECT 244.425 0.3 244.685 8.7 ;
      RECT 244.935 0.3 245.195 8.7 ;
      RECT 247.995 0.17 248.765 0.43 ;
      RECT 247.995 0.17 248.255 8.7 ;
      RECT 248.505 0.17 248.765 8.7 ;
      RECT 249.015 0.18 249.785 0.88 ;
      RECT 249.015 0.18 249.275 8.7 ;
      RECT 249.525 0.18 249.785 8.7 ;
      RECT 245.445 0.52 245.705 8.7 ;
      RECT 246.975 0 247.235 8.7 ;
      RECT 251.41 0.18 252.18 0.88 ;
      RECT 251.41 0.18 251.67 8.7 ;
      RECT 251.92 0.18 252.18 8.7 ;
      RECT 252.43 0.17 253.2 0.43 ;
      RECT 252.43 0.17 252.69 8.7 ;
      RECT 252.94 0.17 253.2 8.7 ;
      RECT 253.45 0.18 254.22 0.88 ;
      RECT 253.45 0.18 253.71 8.7 ;
      RECT 253.96 0.18 254.22 8.7 ;
      RECT 254.47 0.17 255.24 0.43 ;
      RECT 254.47 0.17 254.73 8.7 ;
      RECT 254.98 0.17 255.24 8.7 ;
      RECT 255.49 0.18 256.26 0.88 ;
      RECT 255.49 0.18 255.75 8.7 ;
      RECT 256 0.18 256.26 8.7 ;
      RECT 256.51 0.17 257.28 0.43 ;
      RECT 256.51 0.17 256.77 8.7 ;
      RECT 257.02 0.17 257.28 8.7 ;
      RECT 257.53 0.18 258.3 0.88 ;
      RECT 257.53 0.18 257.79 8.7 ;
      RECT 258.04 0.18 258.3 8.7 ;
      RECT 258.55 0.17 259.32 0.43 ;
      RECT 258.55 0.17 258.81 8.7 ;
      RECT 259.06 0.17 259.32 8.7 ;
      RECT 259.57 0.18 260.34 0.88 ;
      RECT 259.57 0.18 259.83 8.7 ;
      RECT 260.08 0.18 260.34 8.7 ;
      RECT 260.59 0.17 261.36 0.43 ;
      RECT 260.59 0.17 260.85 8.7 ;
      RECT 261.1 0.17 261.36 8.7 ;
      RECT 261.61 0.18 262.38 0.88 ;
      RECT 261.61 0.18 261.87 8.7 ;
      RECT 262.12 0.18 262.38 8.7 ;
      RECT 262.63 0.17 263.4 0.43 ;
      RECT 262.63 0.17 262.89 8.7 ;
      RECT 263.14 0.17 263.4 8.7 ;
      RECT 263.65 0.18 264.42 0.88 ;
      RECT 263.65 0.18 263.91 8.7 ;
      RECT 264.16 0.18 264.42 8.7 ;
      RECT 264.67 0.17 265.44 0.43 ;
      RECT 264.67 0.17 264.93 8.7 ;
      RECT 265.18 0.17 265.44 8.7 ;
      RECT 265.69 0.18 266.46 0.88 ;
      RECT 265.69 0.18 265.95 8.7 ;
      RECT 266.2 0.18 266.46 8.7 ;
      RECT 266.71 0.17 267.48 0.43 ;
      RECT 266.71 0.17 266.97 8.7 ;
      RECT 267.22 0.17 267.48 8.7 ;
      RECT 267.73 0.18 268.5 0.88 ;
      RECT 267.73 0.18 267.99 8.7 ;
      RECT 268.24 0.18 268.5 8.7 ;
      RECT 268.75 0.17 269.52 0.43 ;
      RECT 268.75 0.17 269.01 8.7 ;
      RECT 269.26 0.17 269.52 8.7 ;
      RECT 269.77 0.18 270.54 0.88 ;
      RECT 269.77 0.18 270.03 8.7 ;
      RECT 270.28 0.18 270.54 8.7 ;
      RECT 270.79 0.17 271.56 0.43 ;
      RECT 270.79 0.17 271.05 8.7 ;
      RECT 271.3 0.17 271.56 8.7 ;
      RECT 271.81 0.18 272.58 0.88 ;
      RECT 271.81 0.18 272.07 8.7 ;
      RECT 272.32 0.18 272.58 8.7 ;
      RECT 272.83 0.17 273.6 0.43 ;
      RECT 272.83 0.17 273.09 8.7 ;
      RECT 273.34 0.17 273.6 8.7 ;
      RECT 273.85 0.18 274.62 0.88 ;
      RECT 273.85 0.18 274.11 8.7 ;
      RECT 274.36 0.18 274.62 8.7 ;
      RECT 247.485 0 247.745 8.7 ;
      RECT 274.87 0.17 275.64 0.43 ;
      RECT 274.87 0.17 275.13 8.7 ;
      RECT 275.38 0.17 275.64 8.7 ;
      RECT 250.035 0.3 250.295 8.7 ;
      RECT 250.545 0.3 250.805 8.7 ;
      RECT 275.37 136.13 275.57 136.94 ;
      RECT 276.195 136.21 276.395 136.94 ;
      RECT 276.605 136.21 276.965 136.94 ;
      RECT 276.91 0.52 277.17 4.315 ;
      RECT 277.175 136.21 277.375 136.94 ;
      RECT 277.83 136.21 278.03 136.94 ;
      RECT 278.085 0.52 278.345 2.82 ;
      RECT 278.24 136.21 278.6 136.94 ;
      RECT 278.895 136.21 279.095 136.94 ;
      RECT 279.39 136.21 279.75 136.94 ;
      RECT 280.325 0.18 281.095 0.88 ;
      RECT 280.325 0.18 280.585 12.9 ;
      RECT 280.835 0.18 281.095 12.9 ;
      RECT 279.615 0.52 279.875 2.82 ;
      RECT 279.96 136.21 280.16 136.94 ;
      RECT 281.345 0.155 282.115 0.445 ;
      RECT 281.345 0.155 281.605 13.21 ;
      RECT 281.855 0.155 282.115 13.21 ;
      RECT 280.615 136.21 280.815 136.94 ;
      RECT 281.025 136.21 281.385 136.94 ;
      RECT 281.595 136.21 281.795 136.94 ;
      RECT 282.25 136.21 282.45 136.94 ;
      RECT 282.66 136.21 283.02 136.94 ;
      RECT 283.315 136.21 283.515 136.94 ;
      RECT 283.81 136.21 284.17 136.94 ;
      RECT 284.05 0.52 284.31 14.115 ;
      RECT 284.38 136.21 284.58 136.94 ;
      RECT 284.56 0.52 284.82 13.45 ;
      RECT 285.035 136.21 285.235 136.94 ;
      RECT 285.58 0.155 286.35 0.445 ;
      RECT 285.58 0.155 285.84 8.665 ;
      RECT 286.09 0.155 286.35 8.665 ;
      RECT 285.07 0.52 285.33 11.315 ;
      RECT 285.445 136.21 285.805 136.94 ;
      RECT 286.015 136.21 286.215 136.94 ;
      RECT 286.6 0.52 286.86 9.955 ;
      RECT 286.67 136.21 286.87 136.94 ;
      RECT 287.08 136.21 287.44 136.94 ;
      RECT 287.735 136.21 287.935 136.94 ;
      RECT 288.23 136.21 288.59 136.94 ;
      RECT 288.64 0.3 288.9 8.7 ;
      RECT 288.8 136.21 289 136.94 ;
      RECT 289.455 136.21 289.655 136.94 ;
      RECT 289.15 0.18 289.92 0.88 ;
      RECT 289.865 136.21 290.225 136.94 ;
      RECT 290.435 136.21 290.635 136.94 ;
      RECT 291.09 136.21 291.29 136.94 ;
      RECT 291.345 0.52 291.605 6.28 ;
      RECT 291.5 136.21 291.86 136.94 ;
      RECT 292.155 136.21 292.355 136.94 ;
      RECT 292.72 0.52 292.98 5.57 ;
      RECT 292.65 136.21 293.01 136.94 ;
      RECT 293.22 136.21 293.42 136.94 ;
      RECT 293.23 0.3 293.49 5.235 ;
      RECT 293.74 0.52 294 7.78 ;
      RECT 293.875 136.21 294.075 136.94 ;
      RECT 294.285 136.21 294.645 136.94 ;
      RECT 294.59 0.52 294.85 4.315 ;
      RECT 294.855 136.21 295.055 136.94 ;
      RECT 295.51 136.21 295.71 136.94 ;
      RECT 295.765 0.52 296.025 2.82 ;
      RECT 295.92 136.21 296.28 136.94 ;
      RECT 296.575 136.21 296.775 136.94 ;
      RECT 297.07 136.21 297.43 136.94 ;
      RECT 298.005 0.18 298.775 0.88 ;
      RECT 298.005 0.18 298.265 12.9 ;
      RECT 298.515 0.18 298.775 12.9 ;
      RECT 297.295 0.52 297.555 2.82 ;
      RECT 297.64 136.21 297.84 136.94 ;
      RECT 299.025 0.155 299.795 0.445 ;
      RECT 299.025 0.155 299.285 13.21 ;
      RECT 299.535 0.155 299.795 13.21 ;
      RECT 298.295 136.21 298.495 136.94 ;
      RECT 298.705 136.21 299.065 136.94 ;
      RECT 299.275 136.21 299.475 136.94 ;
      RECT 299.93 136.21 300.13 136.94 ;
      RECT 300.34 136.21 300.7 136.94 ;
      RECT 300.995 136.21 301.195 136.94 ;
      RECT 301.49 136.21 301.85 136.94 ;
      RECT 301.73 0.52 301.99 14.115 ;
      RECT 302.06 136.21 302.26 136.94 ;
      RECT 302.24 0.52 302.5 13.45 ;
      RECT 302.715 136.21 302.915 136.94 ;
      RECT 303.26 0.155 304.03 0.445 ;
      RECT 303.26 0.155 303.52 8.665 ;
      RECT 303.77 0.155 304.03 8.665 ;
      RECT 302.75 0.52 303.01 11.315 ;
      RECT 303.125 136.21 303.485 136.94 ;
      RECT 303.695 136.21 303.895 136.94 ;
      RECT 304.28 0.52 304.54 9.955 ;
      RECT 304.35 136.21 304.55 136.94 ;
      RECT 304.76 136.21 305.12 136.94 ;
      RECT 305.415 136.21 305.615 136.94 ;
      RECT 305.91 136.21 306.27 136.94 ;
      RECT 306.32 0.3 306.58 8.7 ;
      RECT 306.48 136.21 306.68 136.94 ;
      RECT 307.135 136.21 307.335 136.94 ;
      RECT 306.83 0.18 307.6 0.88 ;
      RECT 307.545 136.21 307.905 136.94 ;
      RECT 308.115 136.21 308.315 136.94 ;
      RECT 308.77 136.21 308.97 136.94 ;
      RECT 309.025 0.52 309.285 6.28 ;
      RECT 309.18 136.21 309.54 136.94 ;
      RECT 309.835 136.21 310.035 136.94 ;
      RECT 310.4 0.52 310.66 5.57 ;
      RECT 310.33 136.21 310.69 136.94 ;
      RECT 310.9 136.21 311.1 136.94 ;
      RECT 310.91 0.3 311.17 5.235 ;
      RECT 311.42 0.52 311.68 7.78 ;
      RECT 311.555 136.21 311.755 136.94 ;
      RECT 311.965 136.21 312.325 136.94 ;
      RECT 312.27 0.52 312.53 4.315 ;
      RECT 312.535 136.21 312.735 136.94 ;
      RECT 313.19 136.21 313.39 136.94 ;
      RECT 313.445 0.52 313.705 2.82 ;
      RECT 313.6 136.21 313.96 136.94 ;
      RECT 314.255 136.21 314.455 136.94 ;
      RECT 314.75 136.21 315.11 136.94 ;
      RECT 315.685 0.18 316.455 0.88 ;
      RECT 315.685 0.18 315.945 12.9 ;
      RECT 316.195 0.18 316.455 12.9 ;
      RECT 314.975 0.52 315.235 2.82 ;
      RECT 315.32 136.21 315.52 136.94 ;
      RECT 316.705 0.155 317.475 0.445 ;
      RECT 316.705 0.155 316.965 13.21 ;
      RECT 317.215 0.155 317.475 13.21 ;
      RECT 315.975 136.21 316.175 136.94 ;
      RECT 316.385 136.21 316.745 136.94 ;
      RECT 316.955 136.21 317.155 136.94 ;
      RECT 317.61 136.21 317.81 136.94 ;
      RECT 318.02 136.21 318.38 136.94 ;
      RECT 318.675 136.21 318.875 136.94 ;
      RECT 319.17 136.21 319.53 136.94 ;
      RECT 319.41 0.52 319.67 14.115 ;
      RECT 319.74 136.21 319.94 136.94 ;
      RECT 319.92 0.52 320.18 13.45 ;
      RECT 320.395 136.21 320.595 136.94 ;
      RECT 320.94 0.155 321.71 0.445 ;
      RECT 320.94 0.155 321.2 8.665 ;
      RECT 321.45 0.155 321.71 8.665 ;
      RECT 320.43 0.52 320.69 11.315 ;
      RECT 320.805 136.21 321.165 136.94 ;
      RECT 321.375 136.21 321.575 136.94 ;
      RECT 321.96 0.52 322.22 9.955 ;
      RECT 322.03 136.21 322.23 136.94 ;
      RECT 322.44 136.21 322.8 136.94 ;
      RECT 323.095 136.21 323.295 136.94 ;
      RECT 323.59 136.21 323.95 136.94 ;
      RECT 324 0.3 324.26 8.7 ;
      RECT 324.16 136.21 324.36 136.94 ;
      RECT 324.815 136.21 325.015 136.94 ;
      RECT 324.51 0.18 325.28 0.88 ;
      RECT 325.225 136.21 325.585 136.94 ;
      RECT 325.795 136.21 325.995 136.94 ;
      RECT 326.45 136.21 326.65 136.94 ;
      RECT 326.705 0.52 326.965 6.28 ;
      RECT 326.86 136.21 327.22 136.94 ;
      RECT 327.515 136.21 327.715 136.94 ;
      RECT 328.08 0.52 328.34 5.57 ;
      RECT 328.01 136.21 328.37 136.94 ;
      RECT 328.58 136.21 328.78 136.94 ;
      RECT 328.59 0.3 328.85 5.235 ;
      RECT 329.1 0.52 329.36 7.78 ;
      RECT 329.235 136.21 329.435 136.94 ;
      RECT 329.645 136.21 330.005 136.94 ;
      RECT 329.95 0.52 330.21 4.315 ;
      RECT 330.215 136.21 330.415 136.94 ;
      RECT 330.87 136.21 331.07 136.94 ;
      RECT 331.125 0.52 331.385 2.82 ;
      RECT 331.28 136.21 331.64 136.94 ;
      RECT 331.935 136.21 332.135 136.94 ;
      RECT 332.43 136.21 332.79 136.94 ;
      RECT 333.365 0.18 334.135 0.88 ;
      RECT 333.365 0.18 333.625 12.9 ;
      RECT 333.875 0.18 334.135 12.9 ;
      RECT 332.655 0.52 332.915 2.82 ;
      RECT 333 136.21 333.2 136.94 ;
      RECT 334.385 0.155 335.155 0.445 ;
      RECT 334.385 0.155 334.645 13.21 ;
      RECT 334.895 0.155 335.155 13.21 ;
      RECT 333.655 136.21 333.855 136.94 ;
      RECT 334.065 136.21 334.425 136.94 ;
      RECT 334.635 136.21 334.835 136.94 ;
      RECT 335.29 136.21 335.49 136.94 ;
      RECT 335.7 136.21 336.06 136.94 ;
      RECT 336.355 136.21 336.555 136.94 ;
      RECT 336.85 136.21 337.21 136.94 ;
      RECT 337.09 0.52 337.35 14.115 ;
      RECT 337.42 136.21 337.62 136.94 ;
      RECT 337.6 0.52 337.86 13.45 ;
      RECT 338.075 136.21 338.275 136.94 ;
      RECT 338.62 0.155 339.39 0.445 ;
      RECT 338.62 0.155 338.88 8.665 ;
      RECT 339.13 0.155 339.39 8.665 ;
      RECT 338.11 0.52 338.37 11.315 ;
      RECT 338.485 136.21 338.845 136.94 ;
      RECT 339.055 136.21 339.255 136.94 ;
      RECT 339.64 0.52 339.9 9.955 ;
      RECT 339.71 136.21 339.91 136.94 ;
      RECT 340.12 136.21 340.48 136.94 ;
      RECT 340.775 136.21 340.975 136.94 ;
      RECT 341.27 136.21 341.63 136.94 ;
      RECT 341.68 0.3 341.94 8.7 ;
      RECT 341.84 136.21 342.04 136.94 ;
      RECT 342.495 136.21 342.695 136.94 ;
      RECT 342.19 0.18 342.96 0.88 ;
      RECT 342.905 136.21 343.265 136.94 ;
      RECT 343.475 136.21 343.675 136.94 ;
      RECT 344.13 136.21 344.33 136.94 ;
      RECT 344.385 0.52 344.645 6.28 ;
      RECT 344.54 136.21 344.9 136.94 ;
      RECT 345.195 136.21 345.395 136.94 ;
      RECT 345.76 0.52 346.02 5.57 ;
      RECT 345.69 136.21 346.05 136.94 ;
      RECT 346.26 136.21 346.46 136.94 ;
      RECT 346.27 0.3 346.53 5.235 ;
      RECT 346.78 0.52 347.04 7.78 ;
      RECT 346.915 136.21 347.115 136.94 ;
      RECT 347.325 136.21 347.685 136.94 ;
      RECT 347.63 0.52 347.89 4.315 ;
      RECT 347.895 136.21 348.095 136.94 ;
      RECT 348.55 136.21 348.75 136.94 ;
      RECT 348.805 0.52 349.065 2.82 ;
      RECT 348.96 136.21 349.32 136.94 ;
      RECT 349.615 136.21 349.815 136.94 ;
      RECT 350.11 136.21 350.47 136.94 ;
      RECT 351.045 0.18 351.815 0.88 ;
      RECT 351.045 0.18 351.305 12.9 ;
      RECT 351.555 0.18 351.815 12.9 ;
      RECT 350.335 0.52 350.595 2.82 ;
      RECT 350.68 136.21 350.88 136.94 ;
      RECT 352.065 0.155 352.835 0.445 ;
      RECT 352.065 0.155 352.325 13.21 ;
      RECT 352.575 0.155 352.835 13.21 ;
      RECT 351.335 136.21 351.535 136.94 ;
      RECT 351.745 136.21 352.105 136.94 ;
      RECT 352.315 136.21 352.515 136.94 ;
      RECT 352.97 136.21 353.17 136.94 ;
      RECT 353.38 136.21 353.74 136.94 ;
      RECT 354.035 136.21 354.235 136.94 ;
      RECT 354.53 136.21 354.89 136.94 ;
      RECT 354.77 0.52 355.03 14.115 ;
      RECT 355.1 136.21 355.3 136.94 ;
      RECT 355.28 0.52 355.54 13.45 ;
      RECT 355.755 136.21 355.955 136.94 ;
      RECT 356.3 0.155 357.07 0.445 ;
      RECT 356.3 0.155 356.56 8.665 ;
      RECT 356.81 0.155 357.07 8.665 ;
      RECT 355.79 0.52 356.05 11.315 ;
      RECT 356.165 136.21 356.525 136.94 ;
      RECT 356.735 136.21 356.935 136.94 ;
      RECT 357.32 0.52 357.58 9.955 ;
      RECT 357.39 136.21 357.59 136.94 ;
      RECT 357.8 136.21 358.16 136.94 ;
      RECT 358.455 136.21 358.655 136.94 ;
      RECT 358.95 136.21 359.31 136.94 ;
      RECT 359.36 0.3 359.62 8.7 ;
      RECT 359.52 136.21 359.72 136.94 ;
      RECT 360.175 136.21 360.375 136.94 ;
      RECT 359.87 0.18 360.64 0.88 ;
      RECT 360.585 136.21 360.945 136.94 ;
      RECT 361.155 136.21 361.355 136.94 ;
      RECT 361.81 136.21 362.01 136.94 ;
      RECT 362.065 0.52 362.325 6.28 ;
      RECT 362.22 136.21 362.58 136.94 ;
      RECT 362.875 136.21 363.075 136.94 ;
      RECT 363.44 0.52 363.7 5.57 ;
      RECT 363.37 136.21 363.73 136.94 ;
      RECT 363.94 136.21 364.14 136.94 ;
      RECT 363.95 0.3 364.21 5.235 ;
      RECT 364.46 0.52 364.72 7.78 ;
      RECT 364.595 136.21 364.795 136.94 ;
      RECT 365.005 136.21 365.365 136.94 ;
      RECT 365.31 0.52 365.57 4.315 ;
      RECT 365.575 136.21 365.775 136.94 ;
      RECT 366.23 136.21 366.43 136.94 ;
      RECT 366.485 0.52 366.745 2.82 ;
      RECT 366.64 136.21 367 136.94 ;
      RECT 367.295 136.21 367.495 136.94 ;
      RECT 367.79 136.21 368.15 136.94 ;
      RECT 368.725 0.18 369.495 0.88 ;
      RECT 368.725 0.18 368.985 12.9 ;
      RECT 369.235 0.18 369.495 12.9 ;
      RECT 368.015 0.52 368.275 2.82 ;
      RECT 368.36 136.21 368.56 136.94 ;
      RECT 369.745 0.155 370.515 0.445 ;
      RECT 369.745 0.155 370.005 13.21 ;
      RECT 370.255 0.155 370.515 13.21 ;
      RECT 369.015 136.21 369.215 136.94 ;
      RECT 369.425 136.21 369.785 136.94 ;
      RECT 369.995 136.21 370.195 136.94 ;
      RECT 370.65 136.21 370.85 136.94 ;
      RECT 371.06 136.21 371.42 136.94 ;
      RECT 371.715 136.21 371.915 136.94 ;
      RECT 372.21 136.21 372.57 136.94 ;
      RECT 372.45 0.52 372.71 14.115 ;
      RECT 372.78 136.21 372.98 136.94 ;
      RECT 372.96 0.52 373.22 13.45 ;
      RECT 373.435 136.21 373.635 136.94 ;
      RECT 373.98 0.155 374.75 0.445 ;
      RECT 373.98 0.155 374.24 8.665 ;
      RECT 374.49 0.155 374.75 8.665 ;
      RECT 373.47 0.52 373.73 11.315 ;
      RECT 373.845 136.21 374.205 136.94 ;
      RECT 374.415 136.21 374.615 136.94 ;
      RECT 375 0.52 375.26 9.955 ;
      RECT 375.07 136.21 375.27 136.94 ;
      RECT 375.48 136.21 375.84 136.94 ;
      RECT 376.135 136.21 376.335 136.94 ;
      RECT 376.63 136.21 376.99 136.94 ;
      RECT 377.04 0.3 377.3 8.7 ;
      RECT 377.2 136.21 377.4 136.94 ;
      RECT 377.855 136.21 378.055 136.94 ;
      RECT 377.55 0.18 378.32 0.88 ;
      RECT 378.265 136.21 378.625 136.94 ;
      RECT 378.835 136.21 379.035 136.94 ;
      RECT 379.49 136.21 379.69 136.94 ;
      RECT 379.745 0.52 380.005 6.28 ;
      RECT 379.9 136.21 380.26 136.94 ;
      RECT 380.555 136.21 380.755 136.94 ;
      RECT 381.12 0.52 381.38 5.57 ;
      RECT 381.05 136.21 381.41 136.94 ;
      RECT 381.62 136.21 381.82 136.94 ;
      RECT 381.63 0.3 381.89 5.235 ;
      RECT 382.14 0.52 382.4 7.78 ;
      RECT 382.275 136.21 382.475 136.94 ;
      RECT 382.685 136.21 383.045 136.94 ;
      RECT 382.99 0.52 383.25 4.315 ;
      RECT 383.255 136.21 383.455 136.94 ;
      RECT 383.91 136.21 384.11 136.94 ;
      RECT 384.165 0.52 384.425 2.82 ;
      RECT 384.32 136.21 384.68 136.94 ;
      RECT 384.975 136.21 385.175 136.94 ;
      RECT 385.47 136.21 385.83 136.94 ;
      RECT 386.405 0.18 387.175 0.88 ;
      RECT 386.405 0.18 386.665 12.9 ;
      RECT 386.915 0.18 387.175 12.9 ;
      RECT 385.695 0.52 385.955 2.82 ;
      RECT 386.04 136.21 386.24 136.94 ;
      RECT 387.425 0.155 388.195 0.445 ;
      RECT 387.425 0.155 387.685 13.21 ;
      RECT 387.935 0.155 388.195 13.21 ;
      RECT 386.695 136.21 386.895 136.94 ;
      RECT 387.105 136.21 387.465 136.94 ;
      RECT 387.675 136.21 387.875 136.94 ;
      RECT 388.33 136.21 388.53 136.94 ;
      RECT 388.74 136.21 389.1 136.94 ;
      RECT 389.395 136.21 389.595 136.94 ;
      RECT 389.89 136.21 390.25 136.94 ;
      RECT 390.13 0.52 390.39 14.115 ;
      RECT 390.46 136.21 390.66 136.94 ;
      RECT 390.64 0.52 390.9 13.45 ;
      RECT 391.115 136.21 391.315 136.94 ;
      RECT 391.66 0.155 392.43 0.445 ;
      RECT 391.66 0.155 391.92 8.665 ;
      RECT 392.17 0.155 392.43 8.665 ;
      RECT 391.15 0.52 391.41 11.315 ;
      RECT 391.525 136.21 391.885 136.94 ;
      RECT 392.095 136.21 392.295 136.94 ;
      RECT 392.68 0.52 392.94 9.955 ;
      RECT 392.75 136.21 392.95 136.94 ;
      RECT 393.16 136.21 393.52 136.94 ;
      RECT 393.815 136.21 394.015 136.94 ;
      RECT 394.31 136.21 394.67 136.94 ;
      RECT 394.72 0.3 394.98 8.7 ;
      RECT 394.88 136.21 395.08 136.94 ;
      RECT 395.535 136.21 395.735 136.94 ;
      RECT 395.23 0.18 396 0.88 ;
      RECT 395.945 136.21 396.305 136.94 ;
      RECT 396.515 136.21 396.715 136.94 ;
      RECT 397.17 136.21 397.37 136.94 ;
      RECT 397.425 0.52 397.685 6.28 ;
      RECT 397.58 136.21 397.94 136.94 ;
      RECT 398.235 136.21 398.435 136.94 ;
      RECT 398.8 0.52 399.06 5.57 ;
      RECT 398.73 136.21 399.09 136.94 ;
      RECT 399.3 136.21 399.5 136.94 ;
      RECT 399.31 0.3 399.57 5.235 ;
      RECT 399.82 0.52 400.08 7.78 ;
      RECT 399.955 136.21 400.155 136.94 ;
      RECT 400.365 136.21 400.725 136.94 ;
      RECT 400.67 0.52 400.93 4.315 ;
      RECT 400.935 136.21 401.135 136.94 ;
      RECT 401.59 136.21 401.79 136.94 ;
      RECT 401.845 0.52 402.105 2.82 ;
      RECT 402 136.21 402.36 136.94 ;
      RECT 402.655 136.21 402.855 136.94 ;
      RECT 403.15 136.21 403.51 136.94 ;
      RECT 404.085 0.18 404.855 0.88 ;
      RECT 404.085 0.18 404.345 12.9 ;
      RECT 404.595 0.18 404.855 12.9 ;
      RECT 403.375 0.52 403.635 2.82 ;
      RECT 403.72 136.21 403.92 136.94 ;
      RECT 405.105 0.155 405.875 0.445 ;
      RECT 405.105 0.155 405.365 13.21 ;
      RECT 405.615 0.155 405.875 13.21 ;
      RECT 404.375 136.21 404.575 136.94 ;
      RECT 404.785 136.21 405.145 136.94 ;
      RECT 405.355 136.21 405.555 136.94 ;
      RECT 406.01 136.21 406.21 136.94 ;
      RECT 406.42 136.21 406.78 136.94 ;
      RECT 407.075 136.21 407.275 136.94 ;
      RECT 407.57 136.21 407.93 136.94 ;
      RECT 407.81 0.52 408.07 14.115 ;
      RECT 408.14 136.21 408.34 136.94 ;
      RECT 408.32 0.52 408.58 13.45 ;
      RECT 408.795 136.21 408.995 136.94 ;
      RECT 409.34 0.155 410.11 0.445 ;
      RECT 409.34 0.155 409.6 8.665 ;
      RECT 409.85 0.155 410.11 8.665 ;
      RECT 408.83 0.52 409.09 11.315 ;
      RECT 409.205 136.21 409.565 136.94 ;
      RECT 409.775 136.21 409.975 136.94 ;
      RECT 410.36 0.52 410.62 9.955 ;
      RECT 410.43 136.21 410.63 136.94 ;
      RECT 410.84 136.21 411.2 136.94 ;
      RECT 411.495 136.21 411.695 136.94 ;
      RECT 411.99 136.21 412.35 136.94 ;
      RECT 412.4 0.3 412.66 8.7 ;
      RECT 412.56 136.21 412.76 136.94 ;
      RECT 413.215 136.21 413.415 136.94 ;
      RECT 412.91 0.18 413.68 0.88 ;
      RECT 413.625 136.21 413.985 136.94 ;
      RECT 414.195 136.21 414.395 136.94 ;
      RECT 414.85 136.21 415.05 136.94 ;
      RECT 415.105 0.52 415.365 6.28 ;
      RECT 415.26 136.21 415.62 136.94 ;
      RECT 415.915 136.21 416.115 136.94 ;
      RECT 416.48 0.52 416.74 5.57 ;
      RECT 416.41 136.21 416.77 136.94 ;
      RECT 416.98 136.21 417.18 136.94 ;
      RECT 416.99 0.3 417.25 5.235 ;
      RECT 417.5 0.52 417.76 7.78 ;
      RECT 417.635 136.21 417.835 136.94 ;
      RECT 418.045 136.21 418.405 136.94 ;
      RECT 418.615 136.21 418.815 136.94 ;
      RECT 419.44 53.41 419.64 136.94 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 415.625 0 416.22 136.97 ;
      RECT 416.99 0.3 417.25 136.97 ;
      RECT 418.02 0 419.95 136.97 ;
      RECT 0 0.52 419.95 136.97 ;
      RECT 410.88 0 414.845 136.97 ;
      RECT 409.34 0.155 410.11 136.97 ;
      RECT 403.895 0 407.55 136.97 ;
      RECT 402.365 0 403.115 136.97 ;
      RECT 401.19 0 401.585 136.97 ;
      RECT 399.31 0.3 399.57 136.97 ;
      RECT 397.945 0 398.54 136.97 ;
      RECT 393.2 0 397.165 136.97 ;
      RECT 391.66 0.155 392.43 136.97 ;
      RECT 386.215 0 389.87 136.97 ;
      RECT 384.685 0 385.435 136.97 ;
      RECT 383.51 0 383.905 136.97 ;
      RECT 381.63 0.3 381.89 136.97 ;
      RECT 380.265 0 380.86 136.97 ;
      RECT 375.52 0 379.485 136.97 ;
      RECT 373.98 0.155 374.75 136.97 ;
      RECT 368.535 0 372.19 136.97 ;
      RECT 367.005 0 367.755 136.97 ;
      RECT 365.83 0 366.225 136.97 ;
      RECT 363.95 0.3 364.21 136.97 ;
      RECT 362.585 0 363.18 136.97 ;
      RECT 357.84 0 361.805 136.97 ;
      RECT 356.3 0.155 357.07 136.97 ;
      RECT 350.855 0 354.51 136.97 ;
      RECT 349.325 0 350.075 136.97 ;
      RECT 348.15 0 348.545 136.97 ;
      RECT 346.27 0.3 346.53 136.97 ;
      RECT 344.905 0 345.5 136.97 ;
      RECT 340.16 0 344.125 136.97 ;
      RECT 338.62 0.155 339.39 136.97 ;
      RECT 333.175 0 336.83 136.97 ;
      RECT 331.645 0 332.395 136.97 ;
      RECT 330.47 0 330.865 136.97 ;
      RECT 328.59 0.3 328.85 136.97 ;
      RECT 327.225 0 327.82 136.97 ;
      RECT 322.48 0 326.445 136.97 ;
      RECT 320.94 0.155 321.71 136.97 ;
      RECT 315.495 0 319.15 136.97 ;
      RECT 313.965 0 314.715 136.97 ;
      RECT 312.79 0 313.185 136.97 ;
      RECT 310.91 0.3 311.17 136.97 ;
      RECT 309.545 0 310.14 136.97 ;
      RECT 304.8 0 308.765 136.97 ;
      RECT 303.26 0.155 304.03 136.97 ;
      RECT 297.815 0 301.47 136.97 ;
      RECT 296.285 0 297.035 136.97 ;
      RECT 295.11 0 295.505 136.97 ;
      RECT 293.23 0.3 293.49 136.97 ;
      RECT 291.865 0 292.46 136.97 ;
      RECT 287.12 0 291.085 136.97 ;
      RECT 285.58 0.155 286.35 136.97 ;
      RECT 280.135 0 283.79 136.97 ;
      RECT 278.605 0 279.355 136.97 ;
      RECT 277.43 0 277.825 136.97 ;
      RECT 245.955 0.18 276.65 136.97 ;
      RECT 245.965 0 276.65 136.97 ;
      RECT 238.305 0.3 245.195 136.97 ;
      RECT 232.695 0.3 233.975 136.97 ;
      RECT 230.145 0.3 231.425 136.97 ;
      RECT 228.615 0.3 228.875 136.97 ;
      RECT 225.555 0.3 225.815 136.97 ;
      RECT 224.025 0.3 224.285 136.97 ;
      RECT 215.865 0.3 222.755 136.97 ;
      RECT 206.375 0 213.575 136.97 ;
      RECT 197.195 0.3 204.085 136.97 ;
      RECT 197.205 0 204.085 136.97 ;
      RECT 195.665 0.3 195.925 136.97 ;
      RECT 194.135 0.3 194.395 136.97 ;
      RECT 191.075 0.3 191.335 136.97 ;
      RECT 188.525 0.3 189.805 136.97 ;
      RECT 185.975 0.3 187.255 136.97 ;
      RECT 174.755 0.3 181.645 136.97 ;
      RECT 174.765 0 181.645 136.97 ;
      RECT 143.3 0.18 173.995 136.97 ;
      RECT 142.125 0 142.52 136.97 ;
      RECT 140.595 0 141.345 136.97 ;
      RECT 136.16 0 139.815 136.97 ;
      RECT 133.6 0.155 134.37 136.97 ;
      RECT 128.865 0 132.83 136.97 ;
      RECT 127.49 0 128.085 136.97 ;
      RECT 126.46 0.3 126.72 136.97 ;
      RECT 124.445 0 124.84 136.97 ;
      RECT 122.915 0 123.665 136.97 ;
      RECT 118.48 0 122.135 136.97 ;
      RECT 115.92 0.155 116.69 136.97 ;
      RECT 111.185 0 115.15 136.97 ;
      RECT 109.81 0 110.405 136.97 ;
      RECT 108.78 0.3 109.04 136.97 ;
      RECT 106.765 0 107.16 136.97 ;
      RECT 105.235 0 105.985 136.97 ;
      RECT 100.8 0 104.455 136.97 ;
      RECT 98.24 0.155 99.01 136.97 ;
      RECT 93.505 0 97.47 136.97 ;
      RECT 92.13 0 92.725 136.97 ;
      RECT 91.1 0.3 91.36 136.97 ;
      RECT 89.085 0 89.48 136.97 ;
      RECT 87.555 0 88.305 136.97 ;
      RECT 83.12 0 86.775 136.97 ;
      RECT 80.56 0.155 81.33 136.97 ;
      RECT 75.825 0 79.79 136.97 ;
      RECT 74.45 0 75.045 136.97 ;
      RECT 73.42 0.3 73.68 136.97 ;
      RECT 71.405 0 71.8 136.97 ;
      RECT 69.875 0 70.625 136.97 ;
      RECT 65.44 0 69.095 136.97 ;
      RECT 62.88 0.155 63.65 136.97 ;
      RECT 58.145 0 62.11 136.97 ;
      RECT 56.77 0 57.365 136.97 ;
      RECT 55.74 0.3 56 136.97 ;
      RECT 53.725 0 54.12 136.97 ;
      RECT 52.195 0 52.945 136.97 ;
      RECT 47.76 0 51.415 136.97 ;
      RECT 45.2 0.155 45.97 136.97 ;
      RECT 40.465 0 44.43 136.97 ;
      RECT 39.09 0 39.685 136.97 ;
      RECT 38.06 0.3 38.32 136.97 ;
      RECT 36.045 0 36.44 136.97 ;
      RECT 34.515 0 35.265 136.97 ;
      RECT 30.08 0 33.735 136.97 ;
      RECT 27.52 0.155 28.29 136.97 ;
      RECT 22.785 0 26.75 136.97 ;
      RECT 21.41 0 22.005 136.97 ;
      RECT 20.38 0.3 20.64 136.97 ;
      RECT 18.365 0 18.76 136.97 ;
      RECT 16.835 0 17.585 136.97 ;
      RECT 12.4 0 16.055 136.97 ;
      RECT 9.84 0.155 10.61 136.97 ;
      RECT 5.105 0 9.07 136.97 ;
      RECT 3.73 0 4.325 136.97 ;
      RECT 2.7 0.3 2.96 136.97 ;
      RECT 0 0 1.93 136.97 ;
      RECT 417 0 417.24 136.97 ;
      RECT 399.32 0 399.56 136.97 ;
      RECT 381.64 0 381.88 136.97 ;
      RECT 363.96 0 364.2 136.97 ;
      RECT 346.28 0 346.52 136.97 ;
      RECT 328.6 0 328.84 136.97 ;
      RECT 310.92 0 311.16 136.97 ;
      RECT 293.24 0 293.48 136.97 ;
      RECT 238.305 0 245.185 136.97 ;
      RECT 232.705 0 233.965 136.97 ;
      RECT 230.155 0 231.415 136.97 ;
      RECT 228.625 0 228.865 136.97 ;
      RECT 225.565 0 225.805 136.97 ;
      RECT 224.035 0 224.275 136.97 ;
      RECT 215.865 0 222.745 136.97 ;
      RECT 195.675 0 195.915 136.97 ;
      RECT 194.145 0 194.385 136.97 ;
      RECT 191.085 0 191.325 136.97 ;
      RECT 188.535 0 189.795 136.97 ;
      RECT 185.985 0 187.245 136.97 ;
      RECT 126.47 0 126.71 136.97 ;
      RECT 108.79 0 109.03 136.97 ;
      RECT 91.11 0 91.35 136.97 ;
      RECT 73.43 0 73.67 136.97 ;
      RECT 55.75 0 55.99 136.97 ;
      RECT 38.07 0 38.31 136.97 ;
      RECT 20.39 0 20.63 136.97 ;
      RECT 2.71 0 2.95 136.97 ;
      RECT 143.3 0 173.985 136.97 ;
      RECT 409.35 0 410.1 136.97 ;
      RECT 391.67 0 392.42 136.97 ;
      RECT 373.99 0 374.74 136.97 ;
      RECT 356.31 0 357.06 136.97 ;
      RECT 338.63 0 339.38 136.97 ;
      RECT 320.95 0 321.7 136.97 ;
      RECT 303.27 0 304.02 136.97 ;
      RECT 285.59 0 286.34 136.97 ;
      RECT 133.61 0 134.36 136.97 ;
      RECT 115.93 0 116.68 136.97 ;
      RECT 98.25 0 99 136.97 ;
      RECT 80.57 0 81.32 136.97 ;
      RECT 62.89 0 63.64 136.97 ;
      RECT 45.21 0 45.96 136.97 ;
      RECT 27.53 0 28.28 136.97 ;
      RECT 9.85 0 10.6 136.97 ;
    LAYER Metal3 ;
      RECT 0 0 419.95 136.97 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 250.265 0 276.525 136.97 ;
      RECT 245.115 0 246.935 136.97 ;
      RECT 239.965 0 241.785 136.97 ;
      RECT 414.065 0 419.95 136.97 ;
      RECT 405.225 0 409.125 136.97 ;
      RECT 405.225 47.305 419.95 53.15 ;
      RECT 396.385 0 400.285 136.97 ;
      RECT 387.545 0 391.445 136.97 ;
      RECT 387.545 47.305 400.285 53.15 ;
      RECT 378.705 0 382.605 136.97 ;
      RECT 369.865 0 373.765 136.97 ;
      RECT 369.865 47.305 382.605 53.15 ;
      RECT 361.025 0 364.925 136.97 ;
      RECT 352.185 0 356.085 136.97 ;
      RECT 352.185 47.305 364.925 53.15 ;
      RECT 343.345 0 347.245 136.97 ;
      RECT 334.505 0 338.405 136.97 ;
      RECT 334.505 47.305 347.245 53.15 ;
      RECT 325.665 0 329.565 136.97 ;
      RECT 316.825 0 320.725 136.97 ;
      RECT 316.825 47.305 329.565 53.15 ;
      RECT 307.985 0 311.885 136.97 ;
      RECT 299.145 0 303.045 136.97 ;
      RECT 299.145 47.305 311.885 53.15 ;
      RECT 290.305 0 294.205 136.97 ;
      RECT 281.465 0 285.365 136.97 ;
      RECT 281.465 47.305 294.205 53.15 ;
      RECT 234.815 0 236.635 136.97 ;
      RECT 229.665 0 231.485 136.97 ;
      RECT 224.515 0 226.335 136.97 ;
      RECT 219.365 0 221.185 136.97 ;
      RECT 214.215 0 216.035 136.97 ;
      RECT 209.065 0 210.885 136.97 ;
      RECT 203.915 0 205.735 136.97 ;
      RECT 198.765 0 200.585 136.97 ;
      RECT 193.615 0 195.435 136.97 ;
      RECT 188.465 0 190.285 136.97 ;
      RECT 183.315 0 185.135 136.97 ;
      RECT 178.165 0 179.985 136.97 ;
      RECT 173.015 0 174.835 136.97 ;
      RECT 143.425 0 169.685 136.97 ;
      RECT 134.585 0 138.485 136.97 ;
      RECT 125.745 0 129.645 136.97 ;
      RECT 125.745 47.305 138.485 53.15 ;
      RECT 116.905 0 120.805 136.97 ;
      RECT 108.065 0 111.965 136.97 ;
      RECT 108.065 47.305 120.805 53.15 ;
      RECT 99.225 0 103.125 136.97 ;
      RECT 90.385 0 94.285 136.97 ;
      RECT 90.385 47.305 103.125 53.15 ;
      RECT 81.545 0 85.445 136.97 ;
      RECT 72.705 0 76.605 136.97 ;
      RECT 72.705 47.305 85.445 53.15 ;
      RECT 63.865 0 67.765 136.97 ;
      RECT 55.025 0 58.925 136.97 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 136.97 ;
      RECT 37.345 0 41.245 136.97 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 136.97 ;
      RECT 19.665 0 23.565 136.97 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 136.97 ;
      RECT 0 0 5.885 136.97 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_256x16_c2_bm_bist

END LIBRARY
