# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Thu Aug 21 20:49:12 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_256x32_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_256x32_c2_bm_bist 0 0 ;
  SIZE 416.64 BY 118.78 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 244.49 0 244.75 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171.89 0 172.15 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 243.635 0 243.895 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.745 0 173.005 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 236.65 0 236.91 0.26 ;
    END
  END A_BM[16]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.73 0 179.99 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 238.025 0 238.285 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.355 0 178.615 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 237.16 0 237.42 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.22 0 179.48 0.26 ;
    END
  END A_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 403.95 0 406.76 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.71 0 395.52 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 381.47 0 384.28 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.23 0 373.04 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.99 0 361.8 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.75 0 350.56 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 336.51 0 339.32 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.27 0 328.08 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.03 0 316.84 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.79 0 305.6 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 291.55 0 294.36 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.31 0 283.12 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.07 0 271.88 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 257.83 0 260.64 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.59 0 249.4 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.35 0 238.16 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.94 0 227.75 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.64 0 217.45 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 199.19 0 202 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 188.89 0 191.7 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.48 0 181.29 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.24 0 170.05 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156 0 158.81 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 144.76 0 147.57 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.52 0 136.33 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.28 0 125.09 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.04 0 113.85 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.8 0 102.61 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 118.78 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 0 412.38 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 0 401.14 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 0 389.9 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 0 378.66 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 0 367.42 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 0 356.18 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 0 344.94 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 0 333.7 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 0 322.46 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 0 311.22 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 0 299.98 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 0 288.74 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 0 277.5 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 0 266.26 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 0 255.02 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 0 243.78 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.79 0 222.6 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.49 0 212.3 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 204.34 0 207.15 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 194.04 0 196.85 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 0 175.67 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 0 164.43 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 0 153.19 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 0 141.95 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 0 130.71 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 0 119.47 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 0 108.23 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 0 96.99 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 38.825 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 45.465 412.38 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 45.465 401.14 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 45.465 389.9 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 45.465 378.66 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 45.465 367.42 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 45.465 356.18 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 45.465 344.94 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 45.465 333.7 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 45.465 322.46 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 45.465 311.22 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 45.465 299.98 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 45.465 288.74 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 45.465 277.5 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 45.465 266.26 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 45.465 255.02 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 45.465 243.78 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 45.465 175.67 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 45.465 164.43 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 45.465 153.19 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 45.465 141.95 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 45.465 130.71 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 45.465 119.47 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 45.465 108.23 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 45.465 96.99 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 45.465 85.75 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 45.465 74.51 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 45.465 63.27 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 45.465 52.03 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 45.465 40.79 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 45.465 29.55 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 45.465 18.31 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 45.465 7.07 118.78 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 255.73 0 255.99 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.65 0 160.91 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 254.875 0 255.135 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.505 0 161.765 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 247.89 0 248.15 0.26 ;
    END
  END A_BM[17]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.49 0 168.75 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.265 0 249.525 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.115 0 167.375 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.4 0 248.66 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.98 0 168.24 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.97 0 267.23 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 149.41 0 149.67 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.115 0 266.375 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.265 0 150.525 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.13 0 259.39 0.26 ;
    END
  END A_BM[18]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.25 0 157.51 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 260.505 0 260.765 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.875 0 156.135 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.64 0 259.9 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.74 0 157 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 278.21 0 278.47 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 138.17 0 138.43 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.355 0 277.615 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 139.025 0 139.285 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 270.37 0 270.63 0.26 ;
    END
  END A_BM[19]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.01 0 146.27 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 271.745 0 272.005 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.635 0 144.895 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 270.88 0 271.14 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.5 0 145.76 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 289.45 0 289.71 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.93 0 127.19 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 288.595 0 288.855 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 127.785 0 128.045 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 281.61 0 281.87 0.26 ;
    END
  END A_BM[20]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.77 0 135.03 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.985 0 283.245 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.395 0 133.655 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.12 0 282.38 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.26 0 134.52 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 300.69 0 300.95 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.69 0 115.95 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 299.835 0 300.095 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.545 0 116.805 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 292.85 0 293.11 0.26 ;
    END
  END A_BM[21]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.53 0 123.79 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.225 0 294.485 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.155 0 122.415 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.36 0 293.62 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.02 0 123.28 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.93 0 312.19 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.45 0 104.71 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.075 0 311.335 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 105.305 0 105.565 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.09 0 304.35 0.26 ;
    END
  END A_BM[22]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.29 0 112.55 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 305.465 0 305.725 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.915 0 111.175 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.6 0 304.86 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.78 0 112.04 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 323.17 0 323.43 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 93.21 0 93.47 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 322.315 0 322.575 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 94.065 0 94.325 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.33 0 315.59 0.26 ;
    END
  END A_BM[23]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.05 0 101.31 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 316.705 0 316.965 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.675 0 99.935 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.84 0 316.1 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.54 0 100.8 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.41 0 334.67 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.97 0 82.23 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.555 0 333.815 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.825 0 83.085 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 326.57 0 326.83 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.81 0 90.07 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.945 0 328.205 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.435 0 88.695 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.08 0 327.34 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.3 0 89.56 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 345.65 0 345.91 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.73 0 70.99 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 344.795 0 345.055 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 71.585 0 71.845 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.81 0 338.07 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.57 0 78.83 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.185 0 339.445 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.195 0 77.455 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.32 0 338.58 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.06 0 78.32 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.89 0 357.15 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 59.49 0 59.75 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.035 0 356.295 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.345 0 60.605 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.05 0 349.31 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.33 0 67.59 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 350.425 0 350.685 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 65.955 0 66.215 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.56 0 349.82 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.82 0 67.08 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.13 0 368.39 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 48.25 0 48.51 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 367.275 0 367.535 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 49.105 0 49.365 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.29 0 360.55 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.09 0 56.35 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 361.665 0 361.925 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.715 0 54.975 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.8 0 361.06 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.58 0 55.84 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.37 0 379.63 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.01 0 37.27 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.515 0 378.775 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.865 0 38.125 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.53 0 371.79 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.85 0 45.11 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.905 0 373.165 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 43.475 0 43.735 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.04 0 372.3 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.34 0 44.6 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.61 0 390.87 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 25.77 0 26.03 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 389.755 0 390.015 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 26.625 0 26.885 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.77 0 383.03 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.61 0 33.87 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.145 0 384.405 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.235 0 32.495 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 383.28 0 383.54 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.1 0 33.36 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.85 0 402.11 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.53 0 14.79 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.995 0 401.255 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.385 0 15.645 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.01 0 394.27 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.37 0 22.63 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 395.385 0 395.645 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.995 0 21.255 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.52 0 394.78 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 21.86 0 22.12 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 413.09 0 413.35 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.29 0 3.55 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 412.235 0 412.495 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.145 0 4.405 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.25 0 405.51 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.13 0 11.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 406.625 0 406.885 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.755 0 10.015 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.76 0 406.02 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.62 0 10.88 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 45.223301 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.52 0 204.78 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.184466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 209.11 0 209.37 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 39.656958 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.01 0 204.27 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.618123 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 208.6 0 208.86 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.17 0 212.43 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.68 0 212.94 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.15 0 211.41 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.66 0 211.92 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.63754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.72 0 214.98 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.317152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.21 0 214.47 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 70.245955 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.7 0 213.96 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 68.925566 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.19 0 213.45 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 55.436893 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.28 0 192.54 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 54.065721 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.79 0 193.05 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 62.724919 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.3 0 193.56 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.404531 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.81 0 194.07 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.48 0 202.74 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.796863 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.05 0 206.31 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.54 0 205.8 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.99 0 203.25 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 18.532819 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.41 0 224.67 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 203.31695 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.17 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.213636 LAYER Metal2 ;
      ANTENNAMAXAREACAR 17.755869 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.03 0 205.29 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.95 0 201.21 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.58 0 207.84 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.07 0 207.33 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 201.46 0 201.72 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 416.64 118.78 ;
    LAYER Metal2 ;
      RECT 0.105 45.465 0.305 118.755 ;
      RECT 1.1 118.025 1.3 118.755 ;
      RECT 3.29 0.52 3.55 5.16 ;
      RECT 2.77 4.9 3.55 5.16 ;
      RECT 2.77 4.9 3.03 6.64 ;
      RECT 1.92 118.025 2.12 118.755 ;
      RECT 2.415 118.025 2.615 118.755 ;
      RECT 2.915 118.025 3.115 118.755 ;
      RECT 3.415 118.025 3.615 118.755 ;
      RECT 3.91 118.025 4.11 118.755 ;
      RECT 4.655 0.17 5.425 0.94 ;
      RECT 4.655 0.17 4.915 12.9 ;
      RECT 5.165 0.17 5.425 12.9 ;
      RECT 4.145 0.52 4.405 5.815 ;
      RECT 4.73 118.025 4.93 118.755 ;
      RECT 5.675 0.17 6.445 0.43 ;
      RECT 5.675 0.17 5.935 11.5 ;
      RECT 6.185 0.17 6.445 11.5 ;
      RECT 5.225 118.025 5.425 118.755 ;
      RECT 5.725 118.025 5.925 118.755 ;
      RECT 6.225 118.025 6.425 118.755 ;
      RECT 7.715 0.17 8.485 0.43 ;
      RECT 7.715 0.17 7.975 10.48 ;
      RECT 8.225 0.17 8.485 10.99 ;
      RECT 6.72 118.025 6.92 118.755 ;
      RECT 7.54 118.025 7.74 118.755 ;
      RECT 8.735 0.17 9.505 0.94 ;
      RECT 8.735 0.17 8.995 8.7 ;
      RECT 9.245 0.17 9.505 12.9 ;
      RECT 8.035 118.025 8.235 118.755 ;
      RECT 8.535 118.025 8.735 118.755 ;
      RECT 9.035 118.025 9.235 118.755 ;
      RECT 9.53 118.025 9.73 118.755 ;
      RECT 9.755 0.52 10.015 2.485 ;
      RECT 10.35 118.025 10.55 118.755 ;
      RECT 10.62 0.52 10.88 14.11 ;
      RECT 10.845 118.025 11.045 118.755 ;
      RECT 11.13 0.52 11.39 2.335 ;
      RECT 11.345 118.025 11.545 118.755 ;
      RECT 11.845 118.025 12.045 118.755 ;
      RECT 12.34 118.025 12.54 118.755 ;
      RECT 14.53 0.52 14.79 5.16 ;
      RECT 14.01 4.9 14.79 5.16 ;
      RECT 14.01 4.9 14.27 6.64 ;
      RECT 13.16 118.025 13.36 118.755 ;
      RECT 13.655 118.025 13.855 118.755 ;
      RECT 14.155 118.025 14.355 118.755 ;
      RECT 14.655 118.025 14.855 118.755 ;
      RECT 15.15 118.025 15.35 118.755 ;
      RECT 15.895 0.17 16.665 0.94 ;
      RECT 15.895 0.17 16.155 12.9 ;
      RECT 16.405 0.17 16.665 12.9 ;
      RECT 15.385 0.52 15.645 5.815 ;
      RECT 15.97 118.025 16.17 118.755 ;
      RECT 16.915 0.17 17.685 0.43 ;
      RECT 16.915 0.17 17.175 11.5 ;
      RECT 17.425 0.17 17.685 11.5 ;
      RECT 16.465 118.025 16.665 118.755 ;
      RECT 16.965 118.025 17.165 118.755 ;
      RECT 17.465 118.025 17.665 118.755 ;
      RECT 18.955 0.17 19.725 0.43 ;
      RECT 18.955 0.17 19.215 10.48 ;
      RECT 19.465 0.17 19.725 10.99 ;
      RECT 17.96 118.025 18.16 118.755 ;
      RECT 18.78 118.025 18.98 118.755 ;
      RECT 19.975 0.17 20.745 0.94 ;
      RECT 19.975 0.17 20.235 8.7 ;
      RECT 20.485 0.17 20.745 12.9 ;
      RECT 19.275 118.025 19.475 118.755 ;
      RECT 19.775 118.025 19.975 118.755 ;
      RECT 20.275 118.025 20.475 118.755 ;
      RECT 20.77 118.025 20.97 118.755 ;
      RECT 20.995 0.52 21.255 2.485 ;
      RECT 21.59 118.025 21.79 118.755 ;
      RECT 21.86 0.52 22.12 14.11 ;
      RECT 22.085 118.025 22.285 118.755 ;
      RECT 22.37 0.52 22.63 2.335 ;
      RECT 22.585 118.025 22.785 118.755 ;
      RECT 23.085 118.025 23.285 118.755 ;
      RECT 23.58 118.025 23.78 118.755 ;
      RECT 25.77 0.52 26.03 5.16 ;
      RECT 25.25 4.9 26.03 5.16 ;
      RECT 25.25 4.9 25.51 6.64 ;
      RECT 24.4 118.025 24.6 118.755 ;
      RECT 24.895 118.025 25.095 118.755 ;
      RECT 25.395 118.025 25.595 118.755 ;
      RECT 25.895 118.025 26.095 118.755 ;
      RECT 26.39 118.025 26.59 118.755 ;
      RECT 27.135 0.17 27.905 0.94 ;
      RECT 27.135 0.17 27.395 12.9 ;
      RECT 27.645 0.17 27.905 12.9 ;
      RECT 26.625 0.52 26.885 5.815 ;
      RECT 27.21 118.025 27.41 118.755 ;
      RECT 28.155 0.17 28.925 0.43 ;
      RECT 28.155 0.17 28.415 11.5 ;
      RECT 28.665 0.17 28.925 11.5 ;
      RECT 27.705 118.025 27.905 118.755 ;
      RECT 28.205 118.025 28.405 118.755 ;
      RECT 28.705 118.025 28.905 118.755 ;
      RECT 30.195 0.17 30.965 0.43 ;
      RECT 30.195 0.17 30.455 10.48 ;
      RECT 30.705 0.17 30.965 10.99 ;
      RECT 29.2 118.025 29.4 118.755 ;
      RECT 30.02 118.025 30.22 118.755 ;
      RECT 31.215 0.17 31.985 0.94 ;
      RECT 31.215 0.17 31.475 8.7 ;
      RECT 31.725 0.17 31.985 12.9 ;
      RECT 30.515 118.025 30.715 118.755 ;
      RECT 31.015 118.025 31.215 118.755 ;
      RECT 31.515 118.025 31.715 118.755 ;
      RECT 32.01 118.025 32.21 118.755 ;
      RECT 32.235 0.52 32.495 2.485 ;
      RECT 32.83 118.025 33.03 118.755 ;
      RECT 33.1 0.52 33.36 14.11 ;
      RECT 33.325 118.025 33.525 118.755 ;
      RECT 33.61 0.52 33.87 2.335 ;
      RECT 33.825 118.025 34.025 118.755 ;
      RECT 34.325 118.025 34.525 118.755 ;
      RECT 34.82 118.025 35.02 118.755 ;
      RECT 37.01 0.52 37.27 5.16 ;
      RECT 36.49 4.9 37.27 5.16 ;
      RECT 36.49 4.9 36.75 6.64 ;
      RECT 35.64 118.025 35.84 118.755 ;
      RECT 36.135 118.025 36.335 118.755 ;
      RECT 36.635 118.025 36.835 118.755 ;
      RECT 37.135 118.025 37.335 118.755 ;
      RECT 37.63 118.025 37.83 118.755 ;
      RECT 38.375 0.17 39.145 0.94 ;
      RECT 38.375 0.17 38.635 12.9 ;
      RECT 38.885 0.17 39.145 12.9 ;
      RECT 37.865 0.52 38.125 5.815 ;
      RECT 38.45 118.025 38.65 118.755 ;
      RECT 39.395 0.17 40.165 0.43 ;
      RECT 39.395 0.17 39.655 11.5 ;
      RECT 39.905 0.17 40.165 11.5 ;
      RECT 38.945 118.025 39.145 118.755 ;
      RECT 39.445 118.025 39.645 118.755 ;
      RECT 39.945 118.025 40.145 118.755 ;
      RECT 41.435 0.17 42.205 0.43 ;
      RECT 41.435 0.17 41.695 10.48 ;
      RECT 41.945 0.17 42.205 10.99 ;
      RECT 40.44 118.025 40.64 118.755 ;
      RECT 41.26 118.025 41.46 118.755 ;
      RECT 42.455 0.17 43.225 0.94 ;
      RECT 42.455 0.17 42.715 8.7 ;
      RECT 42.965 0.17 43.225 12.9 ;
      RECT 41.755 118.025 41.955 118.755 ;
      RECT 42.255 118.025 42.455 118.755 ;
      RECT 42.755 118.025 42.955 118.755 ;
      RECT 43.25 118.025 43.45 118.755 ;
      RECT 43.475 0.52 43.735 2.485 ;
      RECT 44.07 118.025 44.27 118.755 ;
      RECT 44.34 0.52 44.6 14.11 ;
      RECT 44.565 118.025 44.765 118.755 ;
      RECT 44.85 0.52 45.11 2.335 ;
      RECT 45.065 118.025 45.265 118.755 ;
      RECT 45.565 118.025 45.765 118.755 ;
      RECT 46.06 118.025 46.26 118.755 ;
      RECT 48.25 0.52 48.51 5.16 ;
      RECT 47.73 4.9 48.51 5.16 ;
      RECT 47.73 4.9 47.99 6.64 ;
      RECT 46.88 118.025 47.08 118.755 ;
      RECT 47.375 118.025 47.575 118.755 ;
      RECT 47.875 118.025 48.075 118.755 ;
      RECT 48.375 118.025 48.575 118.755 ;
      RECT 48.87 118.025 49.07 118.755 ;
      RECT 49.615 0.17 50.385 0.94 ;
      RECT 49.615 0.17 49.875 12.9 ;
      RECT 50.125 0.17 50.385 12.9 ;
      RECT 49.105 0.52 49.365 5.815 ;
      RECT 49.69 118.025 49.89 118.755 ;
      RECT 50.635 0.17 51.405 0.43 ;
      RECT 50.635 0.17 50.895 11.5 ;
      RECT 51.145 0.17 51.405 11.5 ;
      RECT 50.185 118.025 50.385 118.755 ;
      RECT 50.685 118.025 50.885 118.755 ;
      RECT 51.185 118.025 51.385 118.755 ;
      RECT 52.675 0.17 53.445 0.43 ;
      RECT 52.675 0.17 52.935 10.48 ;
      RECT 53.185 0.17 53.445 10.99 ;
      RECT 51.68 118.025 51.88 118.755 ;
      RECT 52.5 118.025 52.7 118.755 ;
      RECT 53.695 0.17 54.465 0.94 ;
      RECT 53.695 0.17 53.955 8.7 ;
      RECT 54.205 0.17 54.465 12.9 ;
      RECT 52.995 118.025 53.195 118.755 ;
      RECT 53.495 118.025 53.695 118.755 ;
      RECT 53.995 118.025 54.195 118.755 ;
      RECT 54.49 118.025 54.69 118.755 ;
      RECT 54.715 0.52 54.975 2.485 ;
      RECT 55.31 118.025 55.51 118.755 ;
      RECT 55.58 0.52 55.84 14.11 ;
      RECT 55.805 118.025 56.005 118.755 ;
      RECT 56.09 0.52 56.35 2.335 ;
      RECT 56.305 118.025 56.505 118.755 ;
      RECT 56.805 118.025 57.005 118.755 ;
      RECT 57.3 118.025 57.5 118.755 ;
      RECT 59.49 0.52 59.75 5.16 ;
      RECT 58.97 4.9 59.75 5.16 ;
      RECT 58.97 4.9 59.23 6.64 ;
      RECT 58.12 118.025 58.32 118.755 ;
      RECT 58.615 118.025 58.815 118.755 ;
      RECT 59.115 118.025 59.315 118.755 ;
      RECT 59.615 118.025 59.815 118.755 ;
      RECT 60.11 118.025 60.31 118.755 ;
      RECT 60.855 0.17 61.625 0.94 ;
      RECT 60.855 0.17 61.115 12.9 ;
      RECT 61.365 0.17 61.625 12.9 ;
      RECT 60.345 0.52 60.605 5.815 ;
      RECT 60.93 118.025 61.13 118.755 ;
      RECT 61.875 0.17 62.645 0.43 ;
      RECT 61.875 0.17 62.135 11.5 ;
      RECT 62.385 0.17 62.645 11.5 ;
      RECT 61.425 118.025 61.625 118.755 ;
      RECT 61.925 118.025 62.125 118.755 ;
      RECT 62.425 118.025 62.625 118.755 ;
      RECT 63.915 0.17 64.685 0.43 ;
      RECT 63.915 0.17 64.175 10.48 ;
      RECT 64.425 0.17 64.685 10.99 ;
      RECT 62.92 118.025 63.12 118.755 ;
      RECT 63.74 118.025 63.94 118.755 ;
      RECT 64.935 0.17 65.705 0.94 ;
      RECT 64.935 0.17 65.195 8.7 ;
      RECT 65.445 0.17 65.705 12.9 ;
      RECT 64.235 118.025 64.435 118.755 ;
      RECT 64.735 118.025 64.935 118.755 ;
      RECT 65.235 118.025 65.435 118.755 ;
      RECT 65.73 118.025 65.93 118.755 ;
      RECT 65.955 0.52 66.215 2.485 ;
      RECT 66.55 118.025 66.75 118.755 ;
      RECT 66.82 0.52 67.08 14.11 ;
      RECT 67.045 118.025 67.245 118.755 ;
      RECT 67.33 0.52 67.59 2.335 ;
      RECT 67.545 118.025 67.745 118.755 ;
      RECT 68.045 118.025 68.245 118.755 ;
      RECT 68.54 118.025 68.74 118.755 ;
      RECT 70.73 0.52 70.99 5.16 ;
      RECT 70.21 4.9 70.99 5.16 ;
      RECT 70.21 4.9 70.47 6.64 ;
      RECT 69.36 118.025 69.56 118.755 ;
      RECT 69.855 118.025 70.055 118.755 ;
      RECT 70.355 118.025 70.555 118.755 ;
      RECT 70.855 118.025 71.055 118.755 ;
      RECT 71.35 118.025 71.55 118.755 ;
      RECT 72.095 0.17 72.865 0.94 ;
      RECT 72.095 0.17 72.355 12.9 ;
      RECT 72.605 0.17 72.865 12.9 ;
      RECT 71.585 0.52 71.845 5.815 ;
      RECT 72.17 118.025 72.37 118.755 ;
      RECT 73.115 0.17 73.885 0.43 ;
      RECT 73.115 0.17 73.375 11.5 ;
      RECT 73.625 0.17 73.885 11.5 ;
      RECT 72.665 118.025 72.865 118.755 ;
      RECT 73.165 118.025 73.365 118.755 ;
      RECT 73.665 118.025 73.865 118.755 ;
      RECT 75.155 0.17 75.925 0.43 ;
      RECT 75.155 0.17 75.415 10.48 ;
      RECT 75.665 0.17 75.925 10.99 ;
      RECT 74.16 118.025 74.36 118.755 ;
      RECT 74.98 118.025 75.18 118.755 ;
      RECT 76.175 0.17 76.945 0.94 ;
      RECT 76.175 0.17 76.435 8.7 ;
      RECT 76.685 0.17 76.945 12.9 ;
      RECT 75.475 118.025 75.675 118.755 ;
      RECT 75.975 118.025 76.175 118.755 ;
      RECT 76.475 118.025 76.675 118.755 ;
      RECT 76.97 118.025 77.17 118.755 ;
      RECT 77.195 0.52 77.455 2.485 ;
      RECT 77.79 118.025 77.99 118.755 ;
      RECT 78.06 0.52 78.32 14.11 ;
      RECT 78.285 118.025 78.485 118.755 ;
      RECT 78.57 0.52 78.83 2.335 ;
      RECT 78.785 118.025 78.985 118.755 ;
      RECT 79.285 118.025 79.485 118.755 ;
      RECT 79.78 118.025 79.98 118.755 ;
      RECT 81.97 0.52 82.23 5.16 ;
      RECT 81.45 4.9 82.23 5.16 ;
      RECT 81.45 4.9 81.71 6.64 ;
      RECT 80.6 118.025 80.8 118.755 ;
      RECT 81.095 118.025 81.295 118.755 ;
      RECT 81.595 118.025 81.795 118.755 ;
      RECT 82.095 118.025 82.295 118.755 ;
      RECT 82.59 118.025 82.79 118.755 ;
      RECT 83.335 0.17 84.105 0.94 ;
      RECT 83.335 0.17 83.595 12.9 ;
      RECT 83.845 0.17 84.105 12.9 ;
      RECT 82.825 0.52 83.085 5.815 ;
      RECT 83.41 118.025 83.61 118.755 ;
      RECT 84.355 0.17 85.125 0.43 ;
      RECT 84.355 0.17 84.615 11.5 ;
      RECT 84.865 0.17 85.125 11.5 ;
      RECT 83.905 118.025 84.105 118.755 ;
      RECT 84.405 118.025 84.605 118.755 ;
      RECT 84.905 118.025 85.105 118.755 ;
      RECT 86.395 0.17 87.165 0.43 ;
      RECT 86.395 0.17 86.655 10.48 ;
      RECT 86.905 0.17 87.165 10.99 ;
      RECT 85.4 118.025 85.6 118.755 ;
      RECT 86.22 118.025 86.42 118.755 ;
      RECT 87.415 0.17 88.185 0.94 ;
      RECT 87.415 0.17 87.675 8.7 ;
      RECT 87.925 0.17 88.185 12.9 ;
      RECT 86.715 118.025 86.915 118.755 ;
      RECT 87.215 118.025 87.415 118.755 ;
      RECT 87.715 118.025 87.915 118.755 ;
      RECT 88.21 118.025 88.41 118.755 ;
      RECT 88.435 0.52 88.695 2.485 ;
      RECT 89.03 118.025 89.23 118.755 ;
      RECT 89.3 0.52 89.56 14.11 ;
      RECT 89.525 118.025 89.725 118.755 ;
      RECT 89.81 0.52 90.07 2.335 ;
      RECT 90.025 118.025 90.225 118.755 ;
      RECT 90.525 118.025 90.725 118.755 ;
      RECT 91.02 118.025 91.22 118.755 ;
      RECT 93.21 0.52 93.47 5.16 ;
      RECT 92.69 4.9 93.47 5.16 ;
      RECT 92.69 4.9 92.95 6.64 ;
      RECT 91.84 118.025 92.04 118.755 ;
      RECT 92.335 118.025 92.535 118.755 ;
      RECT 92.835 118.025 93.035 118.755 ;
      RECT 93.335 118.025 93.535 118.755 ;
      RECT 93.83 118.025 94.03 118.755 ;
      RECT 94.575 0.17 95.345 0.94 ;
      RECT 94.575 0.17 94.835 12.9 ;
      RECT 95.085 0.17 95.345 12.9 ;
      RECT 94.065 0.52 94.325 5.815 ;
      RECT 94.65 118.025 94.85 118.755 ;
      RECT 95.595 0.17 96.365 0.43 ;
      RECT 95.595 0.17 95.855 11.5 ;
      RECT 96.105 0.17 96.365 11.5 ;
      RECT 95.145 118.025 95.345 118.755 ;
      RECT 95.645 118.025 95.845 118.755 ;
      RECT 96.145 118.025 96.345 118.755 ;
      RECT 97.635 0.17 98.405 0.43 ;
      RECT 97.635 0.17 97.895 10.48 ;
      RECT 98.145 0.17 98.405 10.99 ;
      RECT 96.64 118.025 96.84 118.755 ;
      RECT 97.46 118.025 97.66 118.755 ;
      RECT 98.655 0.17 99.425 0.94 ;
      RECT 98.655 0.17 98.915 8.7 ;
      RECT 99.165 0.17 99.425 12.9 ;
      RECT 97.955 118.025 98.155 118.755 ;
      RECT 98.455 118.025 98.655 118.755 ;
      RECT 98.955 118.025 99.155 118.755 ;
      RECT 99.45 118.025 99.65 118.755 ;
      RECT 99.675 0.52 99.935 2.485 ;
      RECT 100.27 118.025 100.47 118.755 ;
      RECT 100.54 0.52 100.8 14.11 ;
      RECT 100.765 118.025 100.965 118.755 ;
      RECT 101.05 0.52 101.31 2.335 ;
      RECT 101.265 118.025 101.465 118.755 ;
      RECT 101.765 118.025 101.965 118.755 ;
      RECT 102.26 118.025 102.46 118.755 ;
      RECT 104.45 0.52 104.71 5.16 ;
      RECT 103.93 4.9 104.71 5.16 ;
      RECT 103.93 4.9 104.19 6.64 ;
      RECT 103.08 118.025 103.28 118.755 ;
      RECT 103.575 118.025 103.775 118.755 ;
      RECT 104.075 118.025 104.275 118.755 ;
      RECT 104.575 118.025 104.775 118.755 ;
      RECT 105.07 118.025 105.27 118.755 ;
      RECT 105.815 0.17 106.585 0.94 ;
      RECT 105.815 0.17 106.075 12.9 ;
      RECT 106.325 0.17 106.585 12.9 ;
      RECT 105.305 0.52 105.565 5.815 ;
      RECT 105.89 118.025 106.09 118.755 ;
      RECT 106.835 0.17 107.605 0.43 ;
      RECT 106.835 0.17 107.095 11.5 ;
      RECT 107.345 0.17 107.605 11.5 ;
      RECT 106.385 118.025 106.585 118.755 ;
      RECT 106.885 118.025 107.085 118.755 ;
      RECT 107.385 118.025 107.585 118.755 ;
      RECT 108.875 0.17 109.645 0.43 ;
      RECT 108.875 0.17 109.135 10.48 ;
      RECT 109.385 0.17 109.645 10.99 ;
      RECT 107.88 118.025 108.08 118.755 ;
      RECT 108.7 118.025 108.9 118.755 ;
      RECT 109.895 0.17 110.665 0.94 ;
      RECT 109.895 0.17 110.155 8.7 ;
      RECT 110.405 0.17 110.665 12.9 ;
      RECT 109.195 118.025 109.395 118.755 ;
      RECT 109.695 118.025 109.895 118.755 ;
      RECT 110.195 118.025 110.395 118.755 ;
      RECT 110.69 118.025 110.89 118.755 ;
      RECT 110.915 0.52 111.175 2.485 ;
      RECT 111.51 118.025 111.71 118.755 ;
      RECT 111.78 0.52 112.04 14.11 ;
      RECT 112.005 118.025 112.205 118.755 ;
      RECT 112.29 0.52 112.55 2.335 ;
      RECT 112.505 118.025 112.705 118.755 ;
      RECT 113.005 118.025 113.205 118.755 ;
      RECT 113.5 118.025 113.7 118.755 ;
      RECT 115.69 0.52 115.95 5.16 ;
      RECT 115.17 4.9 115.95 5.16 ;
      RECT 115.17 4.9 115.43 6.64 ;
      RECT 114.32 118.025 114.52 118.755 ;
      RECT 114.815 118.025 115.015 118.755 ;
      RECT 115.315 118.025 115.515 118.755 ;
      RECT 115.815 118.025 116.015 118.755 ;
      RECT 116.31 118.025 116.51 118.755 ;
      RECT 117.055 0.17 117.825 0.94 ;
      RECT 117.055 0.17 117.315 12.9 ;
      RECT 117.565 0.17 117.825 12.9 ;
      RECT 116.545 0.52 116.805 5.815 ;
      RECT 117.13 118.025 117.33 118.755 ;
      RECT 118.075 0.17 118.845 0.43 ;
      RECT 118.075 0.17 118.335 11.5 ;
      RECT 118.585 0.17 118.845 11.5 ;
      RECT 117.625 118.025 117.825 118.755 ;
      RECT 118.125 118.025 118.325 118.755 ;
      RECT 118.625 118.025 118.825 118.755 ;
      RECT 120.115 0.17 120.885 0.43 ;
      RECT 120.115 0.17 120.375 10.48 ;
      RECT 120.625 0.17 120.885 10.99 ;
      RECT 119.12 118.025 119.32 118.755 ;
      RECT 119.94 118.025 120.14 118.755 ;
      RECT 121.135 0.17 121.905 0.94 ;
      RECT 121.135 0.17 121.395 8.7 ;
      RECT 121.645 0.17 121.905 12.9 ;
      RECT 120.435 118.025 120.635 118.755 ;
      RECT 120.935 118.025 121.135 118.755 ;
      RECT 121.435 118.025 121.635 118.755 ;
      RECT 121.93 118.025 122.13 118.755 ;
      RECT 122.155 0.52 122.415 2.485 ;
      RECT 122.75 118.025 122.95 118.755 ;
      RECT 123.02 0.52 123.28 14.11 ;
      RECT 123.245 118.025 123.445 118.755 ;
      RECT 123.53 0.52 123.79 2.335 ;
      RECT 123.745 118.025 123.945 118.755 ;
      RECT 124.245 118.025 124.445 118.755 ;
      RECT 124.74 118.025 124.94 118.755 ;
      RECT 126.93 0.52 127.19 5.16 ;
      RECT 126.41 4.9 127.19 5.16 ;
      RECT 126.41 4.9 126.67 6.64 ;
      RECT 125.56 118.025 125.76 118.755 ;
      RECT 126.055 118.025 126.255 118.755 ;
      RECT 126.555 118.025 126.755 118.755 ;
      RECT 127.055 118.025 127.255 118.755 ;
      RECT 127.55 118.025 127.75 118.755 ;
      RECT 128.295 0.17 129.065 0.94 ;
      RECT 128.295 0.17 128.555 12.9 ;
      RECT 128.805 0.17 129.065 12.9 ;
      RECT 127.785 0.52 128.045 5.815 ;
      RECT 128.37 118.025 128.57 118.755 ;
      RECT 129.315 0.17 130.085 0.43 ;
      RECT 129.315 0.17 129.575 11.5 ;
      RECT 129.825 0.17 130.085 11.5 ;
      RECT 128.865 118.025 129.065 118.755 ;
      RECT 129.365 118.025 129.565 118.755 ;
      RECT 129.865 118.025 130.065 118.755 ;
      RECT 131.355 0.17 132.125 0.43 ;
      RECT 131.355 0.17 131.615 10.48 ;
      RECT 131.865 0.17 132.125 10.99 ;
      RECT 130.36 118.025 130.56 118.755 ;
      RECT 131.18 118.025 131.38 118.755 ;
      RECT 132.375 0.17 133.145 0.94 ;
      RECT 132.375 0.17 132.635 8.7 ;
      RECT 132.885 0.17 133.145 12.9 ;
      RECT 131.675 118.025 131.875 118.755 ;
      RECT 132.175 118.025 132.375 118.755 ;
      RECT 132.675 118.025 132.875 118.755 ;
      RECT 133.17 118.025 133.37 118.755 ;
      RECT 133.395 0.52 133.655 2.485 ;
      RECT 133.99 118.025 134.19 118.755 ;
      RECT 134.26 0.52 134.52 14.11 ;
      RECT 134.485 118.025 134.685 118.755 ;
      RECT 134.77 0.52 135.03 2.335 ;
      RECT 134.985 118.025 135.185 118.755 ;
      RECT 135.485 118.025 135.685 118.755 ;
      RECT 135.98 118.025 136.18 118.755 ;
      RECT 138.17 0.52 138.43 5.16 ;
      RECT 137.65 4.9 138.43 5.16 ;
      RECT 137.65 4.9 137.91 6.64 ;
      RECT 136.8 118.025 137 118.755 ;
      RECT 137.295 118.025 137.495 118.755 ;
      RECT 137.795 118.025 137.995 118.755 ;
      RECT 138.295 118.025 138.495 118.755 ;
      RECT 138.79 118.025 138.99 118.755 ;
      RECT 139.535 0.17 140.305 0.94 ;
      RECT 139.535 0.17 139.795 12.9 ;
      RECT 140.045 0.17 140.305 12.9 ;
      RECT 139.025 0.52 139.285 5.815 ;
      RECT 139.61 118.025 139.81 118.755 ;
      RECT 140.555 0.17 141.325 0.43 ;
      RECT 140.555 0.17 140.815 11.5 ;
      RECT 141.065 0.17 141.325 11.5 ;
      RECT 140.105 118.025 140.305 118.755 ;
      RECT 140.605 118.025 140.805 118.755 ;
      RECT 141.105 118.025 141.305 118.755 ;
      RECT 142.595 0.17 143.365 0.43 ;
      RECT 142.595 0.17 142.855 10.48 ;
      RECT 143.105 0.17 143.365 10.99 ;
      RECT 141.6 118.025 141.8 118.755 ;
      RECT 142.42 118.025 142.62 118.755 ;
      RECT 143.615 0.17 144.385 0.94 ;
      RECT 143.615 0.17 143.875 8.7 ;
      RECT 144.125 0.17 144.385 12.9 ;
      RECT 142.915 118.025 143.115 118.755 ;
      RECT 143.415 118.025 143.615 118.755 ;
      RECT 143.915 118.025 144.115 118.755 ;
      RECT 144.41 118.025 144.61 118.755 ;
      RECT 144.635 0.52 144.895 2.485 ;
      RECT 145.23 118.025 145.43 118.755 ;
      RECT 145.5 0.52 145.76 14.11 ;
      RECT 145.725 118.025 145.925 118.755 ;
      RECT 146.01 0.52 146.27 2.335 ;
      RECT 146.225 118.025 146.425 118.755 ;
      RECT 146.725 118.025 146.925 118.755 ;
      RECT 147.22 118.025 147.42 118.755 ;
      RECT 149.41 0.52 149.67 5.16 ;
      RECT 148.89 4.9 149.67 5.16 ;
      RECT 148.89 4.9 149.15 6.64 ;
      RECT 148.04 118.025 148.24 118.755 ;
      RECT 148.535 118.025 148.735 118.755 ;
      RECT 149.035 118.025 149.235 118.755 ;
      RECT 149.535 118.025 149.735 118.755 ;
      RECT 150.03 118.025 150.23 118.755 ;
      RECT 150.775 0.17 151.545 0.94 ;
      RECT 150.775 0.17 151.035 12.9 ;
      RECT 151.285 0.17 151.545 12.9 ;
      RECT 150.265 0.52 150.525 5.815 ;
      RECT 150.85 118.025 151.05 118.755 ;
      RECT 151.795 0.17 152.565 0.43 ;
      RECT 151.795 0.17 152.055 11.5 ;
      RECT 152.305 0.17 152.565 11.5 ;
      RECT 151.345 118.025 151.545 118.755 ;
      RECT 151.845 118.025 152.045 118.755 ;
      RECT 152.345 118.025 152.545 118.755 ;
      RECT 153.835 0.17 154.605 0.43 ;
      RECT 153.835 0.17 154.095 10.48 ;
      RECT 154.345 0.17 154.605 10.99 ;
      RECT 152.84 118.025 153.04 118.755 ;
      RECT 153.66 118.025 153.86 118.755 ;
      RECT 154.855 0.17 155.625 0.94 ;
      RECT 154.855 0.17 155.115 8.7 ;
      RECT 155.365 0.17 155.625 12.9 ;
      RECT 154.155 118.025 154.355 118.755 ;
      RECT 154.655 118.025 154.855 118.755 ;
      RECT 155.155 118.025 155.355 118.755 ;
      RECT 155.65 118.025 155.85 118.755 ;
      RECT 155.875 0.52 156.135 2.485 ;
      RECT 156.47 118.025 156.67 118.755 ;
      RECT 156.74 0.52 157 14.11 ;
      RECT 156.965 118.025 157.165 118.755 ;
      RECT 157.25 0.52 157.51 2.335 ;
      RECT 157.465 118.025 157.665 118.755 ;
      RECT 157.965 118.025 158.165 118.755 ;
      RECT 158.46 118.025 158.66 118.755 ;
      RECT 160.65 0.52 160.91 5.16 ;
      RECT 160.13 4.9 160.91 5.16 ;
      RECT 160.13 4.9 160.39 6.64 ;
      RECT 159.28 118.025 159.48 118.755 ;
      RECT 159.775 118.025 159.975 118.755 ;
      RECT 160.275 118.025 160.475 118.755 ;
      RECT 160.775 118.025 160.975 118.755 ;
      RECT 161.27 118.025 161.47 118.755 ;
      RECT 162.015 0.17 162.785 0.94 ;
      RECT 162.015 0.17 162.275 12.9 ;
      RECT 162.525 0.17 162.785 12.9 ;
      RECT 161.505 0.52 161.765 5.815 ;
      RECT 162.09 118.025 162.29 118.755 ;
      RECT 163.035 0.17 163.805 0.43 ;
      RECT 163.035 0.17 163.295 11.5 ;
      RECT 163.545 0.17 163.805 11.5 ;
      RECT 162.585 118.025 162.785 118.755 ;
      RECT 163.085 118.025 163.285 118.755 ;
      RECT 163.585 118.025 163.785 118.755 ;
      RECT 165.075 0.17 165.845 0.43 ;
      RECT 165.075 0.17 165.335 10.48 ;
      RECT 165.585 0.17 165.845 10.99 ;
      RECT 164.08 118.025 164.28 118.755 ;
      RECT 164.9 118.025 165.1 118.755 ;
      RECT 166.095 0.17 166.865 0.94 ;
      RECT 166.095 0.17 166.355 8.7 ;
      RECT 166.605 0.17 166.865 12.9 ;
      RECT 165.395 118.025 165.595 118.755 ;
      RECT 165.895 118.025 166.095 118.755 ;
      RECT 166.395 118.025 166.595 118.755 ;
      RECT 166.89 118.025 167.09 118.755 ;
      RECT 167.115 0.52 167.375 2.485 ;
      RECT 167.71 118.025 167.91 118.755 ;
      RECT 167.98 0.52 168.24 14.11 ;
      RECT 168.205 118.025 168.405 118.755 ;
      RECT 168.49 0.52 168.75 2.335 ;
      RECT 168.705 118.025 168.905 118.755 ;
      RECT 169.205 118.025 169.405 118.755 ;
      RECT 169.7 118.025 169.9 118.755 ;
      RECT 171.89 0.52 172.15 5.16 ;
      RECT 171.37 4.9 172.15 5.16 ;
      RECT 171.37 4.9 171.63 6.64 ;
      RECT 170.52 118.025 170.72 118.755 ;
      RECT 171.015 118.025 171.215 118.755 ;
      RECT 171.515 118.025 171.715 118.755 ;
      RECT 172.015 118.025 172.215 118.755 ;
      RECT 172.51 118.025 172.71 118.755 ;
      RECT 173.255 0.17 174.025 0.94 ;
      RECT 173.255 0.17 173.515 12.9 ;
      RECT 173.765 0.17 174.025 12.9 ;
      RECT 172.745 0.52 173.005 5.815 ;
      RECT 173.33 118.025 173.53 118.755 ;
      RECT 174.275 0.17 175.045 0.43 ;
      RECT 174.275 0.17 174.535 11.5 ;
      RECT 174.785 0.17 175.045 11.5 ;
      RECT 173.825 118.025 174.025 118.755 ;
      RECT 174.325 118.025 174.525 118.755 ;
      RECT 174.825 118.025 175.025 118.755 ;
      RECT 176.315 0.17 177.085 0.43 ;
      RECT 176.315 0.17 176.575 10.48 ;
      RECT 176.825 0.17 177.085 10.99 ;
      RECT 175.32 118.025 175.52 118.755 ;
      RECT 176.14 118.025 176.34 118.755 ;
      RECT 177.335 0.17 178.105 0.94 ;
      RECT 177.335 0.17 177.595 8.7 ;
      RECT 177.845 0.17 178.105 12.9 ;
      RECT 176.635 118.025 176.835 118.755 ;
      RECT 177.135 118.025 177.335 118.755 ;
      RECT 177.635 118.025 177.835 118.755 ;
      RECT 178.13 118.025 178.33 118.755 ;
      RECT 178.355 0.52 178.615 2.485 ;
      RECT 178.95 118.025 179.15 118.755 ;
      RECT 179.22 0.52 179.48 14.11 ;
      RECT 179.445 118.025 179.645 118.755 ;
      RECT 179.73 0.52 179.99 2.335 ;
      RECT 179.945 118.025 180.145 118.755 ;
      RECT 180.445 118.025 180.645 118.755 ;
      RECT 182.435 0.17 183.205 0.43 ;
      RECT 182.435 0.17 182.695 8.7 ;
      RECT 182.945 0.17 183.205 8.7 ;
      RECT 183.455 0.17 184.225 0.94 ;
      RECT 183.455 0.17 183.715 8.7 ;
      RECT 183.965 0.17 184.225 8.7 ;
      RECT 184.475 0.17 185.245 0.43 ;
      RECT 184.475 0.17 184.735 8.7 ;
      RECT 184.985 0.17 185.245 8.7 ;
      RECT 185.495 0.17 186.265 0.94 ;
      RECT 185.495 0.17 185.755 8.7 ;
      RECT 186.005 0.17 186.265 8.7 ;
      RECT 186.515 0.17 187.285 0.43 ;
      RECT 186.515 0.17 186.775 8.7 ;
      RECT 187.025 0.17 187.285 8.7 ;
      RECT 187.535 0.17 188.305 0.94 ;
      RECT 187.535 0.17 187.795 8.7 ;
      RECT 188.045 0.17 188.305 8.7 ;
      RECT 180.94 118.025 181.14 118.755 ;
      RECT 181.76 118.025 181.96 118.755 ;
      RECT 182.755 118.025 182.955 118.755 ;
      RECT 190.24 0.17 191.01 0.94 ;
      RECT 190.24 0.17 190.5 8.7 ;
      RECT 190.75 0.17 191.01 8.7 ;
      RECT 188.71 0.3 188.97 8.7 ;
      RECT 189.22 0 189.48 8.7 ;
      RECT 189.73 0 189.99 8.7 ;
      RECT 191.26 0 191.52 8.7 ;
      RECT 191.77 0 192.03 8.7 ;
      RECT 192.28 0.52 192.54 8.7 ;
      RECT 192.79 0.52 193.05 8.7 ;
      RECT 193.3 0.52 193.56 8.7 ;
      RECT 195.34 0.17 196.11 0.94 ;
      RECT 195.34 0.17 195.6 8.7 ;
      RECT 195.85 0.17 196.11 8.7 ;
      RECT 196.36 0.17 197.13 0.43 ;
      RECT 196.36 0.17 196.62 8.7 ;
      RECT 196.87 0.17 197.13 8.7 ;
      RECT 193.81 0.52 194.07 8.7 ;
      RECT 194.32 0 194.58 8.7 ;
      RECT 194.83 0 195.09 8.7 ;
      RECT 197.38 0.3 197.64 8.7 ;
      RECT 197.89 0.3 198.15 8.7 ;
      RECT 199.93 0.17 200.7 0.94 ;
      RECT 199.93 0.17 200.19 8.7 ;
      RECT 200.44 0.17 200.7 8.7 ;
      RECT 198.4 0.3 198.66 8.7 ;
      RECT 198.91 0.3 199.17 8.7 ;
      RECT 199.42 0.3 199.68 8.7 ;
      RECT 200.95 0.52 201.21 8.7 ;
      RECT 201.46 0.52 201.72 8.7 ;
      RECT 201.97 0.3 202.23 8.7 ;
      RECT 202.48 0.52 202.74 8.7 ;
      RECT 202.99 0.52 203.25 8.7 ;
      RECT 203.5 0.3 203.76 8.7 ;
      RECT 204.01 0.52 204.27 8.7 ;
      RECT 204.52 0.52 204.78 8.7 ;
      RECT 205.03 0.52 205.29 8.7 ;
      RECT 205.54 0.52 205.8 8.7 ;
      RECT 206.05 0.52 206.31 8.7 ;
      RECT 206.56 0.3 206.82 8.7 ;
      RECT 207.07 0.52 207.33 8.7 ;
      RECT 207.58 0.52 207.84 8.7 ;
      RECT 208.09 0.3 208.35 8.7 ;
      RECT 210.13 0.17 210.9 0.94 ;
      RECT 210.13 0.17 210.39 8.7 ;
      RECT 210.64 0.17 210.9 8.7 ;
      RECT 208.6 0.52 208.86 8.7 ;
      RECT 209.11 0.52 209.37 8.7 ;
      RECT 209.62 0.3 209.88 8.7 ;
      RECT 211.15 0.52 211.41 8.7 ;
      RECT 211.66 0.52 211.92 8.7 ;
      RECT 212.17 0.52 212.43 8.7 ;
      RECT 212.68 0.52 212.94 8.7 ;
      RECT 213.19 0.52 213.45 8.7 ;
      RECT 213.7 0.52 213.96 8.7 ;
      RECT 214.21 0.52 214.47 8.7 ;
      RECT 216.25 0.17 217.02 0.94 ;
      RECT 216.25 0.17 216.51 8.7 ;
      RECT 216.76 0.17 217.02 8.7 ;
      RECT 214.72 0.52 214.98 8.7 ;
      RECT 215.23 0 215.49 8.7 ;
      RECT 215.74 0 216 8.7 ;
      RECT 217.27 0 217.53 8.7 ;
      RECT 219.31 0.17 220.08 0.43 ;
      RECT 219.31 0.17 219.57 8.7 ;
      RECT 219.82 0.17 220.08 8.7 ;
      RECT 217.78 0 218.04 8.7 ;
      RECT 218.29 0.3 218.55 8.7 ;
      RECT 218.8 0.3 219.06 8.7 ;
      RECT 220.33 0.3 220.59 8.7 ;
      RECT 220.84 0.3 221.1 8.7 ;
      RECT 221.35 0.3 221.61 8.7 ;
      RECT 221.86 0.3 222.12 8.7 ;
      RECT 222.37 0 222.63 8.7 ;
      RECT 222.88 0 223.14 8.7 ;
      RECT 224.92 0.17 225.69 0.43 ;
      RECT 224.92 0.17 225.18 8.7 ;
      RECT 225.43 0.17 225.69 8.7 ;
      RECT 225.94 0.17 226.71 0.94 ;
      RECT 225.94 0.17 226.2 25.5 ;
      RECT 226.45 0.17 226.71 33.9 ;
      RECT 226.96 0.17 227.73 0.43 ;
      RECT 226.96 0.17 227.22 8.7 ;
      RECT 227.47 0.17 227.73 8.7 ;
      RECT 228.335 0.17 229.105 0.94 ;
      RECT 228.335 0.17 228.595 8.7 ;
      RECT 228.845 0.17 229.105 8.7 ;
      RECT 229.355 0.17 230.125 0.43 ;
      RECT 229.355 0.17 229.615 8.7 ;
      RECT 229.865 0.17 230.125 8.7 ;
      RECT 230.375 0.17 231.145 0.94 ;
      RECT 230.375 0.17 230.635 8.7 ;
      RECT 230.885 0.17 231.145 8.7 ;
      RECT 231.395 0.17 232.165 0.43 ;
      RECT 231.395 0.17 231.655 8.7 ;
      RECT 231.905 0.17 232.165 8.7 ;
      RECT 232.415 0.17 233.185 0.94 ;
      RECT 232.415 0.17 232.675 8.7 ;
      RECT 232.925 0.17 233.185 8.7 ;
      RECT 223.39 0.3 223.65 8.7 ;
      RECT 233.435 0.17 234.205 0.43 ;
      RECT 233.435 0.17 233.695 8.7 ;
      RECT 233.945 0.17 234.205 8.7 ;
      RECT 223.9 0.3 224.16 8.7 ;
      RECT 224.41 0.52 224.67 8.7 ;
      RECT 233.685 118.025 233.885 118.755 ;
      RECT 234.68 118.025 234.88 118.755 ;
      RECT 235.5 118.025 235.7 118.755 ;
      RECT 235.995 118.025 236.195 118.755 ;
      RECT 236.495 118.025 236.695 118.755 ;
      RECT 236.65 0.52 236.91 2.335 ;
      RECT 236.995 118.025 237.195 118.755 ;
      RECT 237.16 0.52 237.42 14.11 ;
      RECT 237.49 118.025 237.69 118.755 ;
      RECT 238.535 0.17 239.305 0.94 ;
      RECT 239.045 0.17 239.305 8.7 ;
      RECT 238.535 0.17 238.795 12.9 ;
      RECT 238.025 0.52 238.285 2.485 ;
      RECT 238.31 118.025 238.51 118.755 ;
      RECT 239.555 0.17 240.325 0.43 ;
      RECT 240.065 0.17 240.325 10.48 ;
      RECT 239.555 0.17 239.815 10.99 ;
      RECT 238.805 118.025 239.005 118.755 ;
      RECT 239.305 118.025 239.505 118.755 ;
      RECT 239.805 118.025 240.005 118.755 ;
      RECT 240.3 118.025 240.5 118.755 ;
      RECT 241.595 0.17 242.365 0.43 ;
      RECT 241.595 0.17 241.855 11.5 ;
      RECT 242.105 0.17 242.365 11.5 ;
      RECT 241.12 118.025 241.32 118.755 ;
      RECT 241.615 118.025 241.815 118.755 ;
      RECT 242.615 0.17 243.385 0.94 ;
      RECT 242.615 0.17 242.875 12.9 ;
      RECT 243.125 0.17 243.385 12.9 ;
      RECT 242.115 118.025 242.315 118.755 ;
      RECT 242.615 118.025 242.815 118.755 ;
      RECT 243.11 118.025 243.31 118.755 ;
      RECT 243.635 0.52 243.895 5.815 ;
      RECT 244.49 0.52 244.75 5.16 ;
      RECT 244.49 4.9 245.27 5.16 ;
      RECT 245.01 4.9 245.27 6.64 ;
      RECT 243.93 118.025 244.13 118.755 ;
      RECT 244.425 118.025 244.625 118.755 ;
      RECT 244.925 118.025 245.125 118.755 ;
      RECT 245.425 118.025 245.625 118.755 ;
      RECT 245.92 118.025 246.12 118.755 ;
      RECT 246.74 118.025 246.94 118.755 ;
      RECT 247.235 118.025 247.435 118.755 ;
      RECT 247.735 118.025 247.935 118.755 ;
      RECT 247.89 0.52 248.15 2.335 ;
      RECT 248.235 118.025 248.435 118.755 ;
      RECT 248.4 0.52 248.66 14.11 ;
      RECT 248.73 118.025 248.93 118.755 ;
      RECT 249.775 0.17 250.545 0.94 ;
      RECT 250.285 0.17 250.545 8.7 ;
      RECT 249.775 0.17 250.035 12.9 ;
      RECT 249.265 0.52 249.525 2.485 ;
      RECT 249.55 118.025 249.75 118.755 ;
      RECT 250.795 0.17 251.565 0.43 ;
      RECT 251.305 0.17 251.565 10.48 ;
      RECT 250.795 0.17 251.055 10.99 ;
      RECT 250.045 118.025 250.245 118.755 ;
      RECT 250.545 118.025 250.745 118.755 ;
      RECT 251.045 118.025 251.245 118.755 ;
      RECT 251.54 118.025 251.74 118.755 ;
      RECT 252.835 0.17 253.605 0.43 ;
      RECT 252.835 0.17 253.095 11.5 ;
      RECT 253.345 0.17 253.605 11.5 ;
      RECT 252.36 118.025 252.56 118.755 ;
      RECT 252.855 118.025 253.055 118.755 ;
      RECT 253.855 0.17 254.625 0.94 ;
      RECT 253.855 0.17 254.115 12.9 ;
      RECT 254.365 0.17 254.625 12.9 ;
      RECT 253.355 118.025 253.555 118.755 ;
      RECT 253.855 118.025 254.055 118.755 ;
      RECT 254.35 118.025 254.55 118.755 ;
      RECT 254.875 0.52 255.135 5.815 ;
      RECT 255.73 0.52 255.99 5.16 ;
      RECT 255.73 4.9 256.51 5.16 ;
      RECT 256.25 4.9 256.51 6.64 ;
      RECT 255.17 118.025 255.37 118.755 ;
      RECT 255.665 118.025 255.865 118.755 ;
      RECT 256.165 118.025 256.365 118.755 ;
      RECT 256.665 118.025 256.865 118.755 ;
      RECT 257.16 118.025 257.36 118.755 ;
      RECT 257.98 118.025 258.18 118.755 ;
      RECT 258.475 118.025 258.675 118.755 ;
      RECT 258.975 118.025 259.175 118.755 ;
      RECT 259.13 0.52 259.39 2.335 ;
      RECT 259.475 118.025 259.675 118.755 ;
      RECT 259.64 0.52 259.9 14.11 ;
      RECT 259.97 118.025 260.17 118.755 ;
      RECT 261.015 0.17 261.785 0.94 ;
      RECT 261.525 0.17 261.785 8.7 ;
      RECT 261.015 0.17 261.275 12.9 ;
      RECT 260.505 0.52 260.765 2.485 ;
      RECT 260.79 118.025 260.99 118.755 ;
      RECT 262.035 0.17 262.805 0.43 ;
      RECT 262.545 0.17 262.805 10.48 ;
      RECT 262.035 0.17 262.295 10.99 ;
      RECT 261.285 118.025 261.485 118.755 ;
      RECT 261.785 118.025 261.985 118.755 ;
      RECT 262.285 118.025 262.485 118.755 ;
      RECT 262.78 118.025 262.98 118.755 ;
      RECT 264.075 0.17 264.845 0.43 ;
      RECT 264.075 0.17 264.335 11.5 ;
      RECT 264.585 0.17 264.845 11.5 ;
      RECT 263.6 118.025 263.8 118.755 ;
      RECT 264.095 118.025 264.295 118.755 ;
      RECT 265.095 0.17 265.865 0.94 ;
      RECT 265.095 0.17 265.355 12.9 ;
      RECT 265.605 0.17 265.865 12.9 ;
      RECT 264.595 118.025 264.795 118.755 ;
      RECT 265.095 118.025 265.295 118.755 ;
      RECT 265.59 118.025 265.79 118.755 ;
      RECT 266.115 0.52 266.375 5.815 ;
      RECT 266.97 0.52 267.23 5.16 ;
      RECT 266.97 4.9 267.75 5.16 ;
      RECT 267.49 4.9 267.75 6.64 ;
      RECT 266.41 118.025 266.61 118.755 ;
      RECT 266.905 118.025 267.105 118.755 ;
      RECT 267.405 118.025 267.605 118.755 ;
      RECT 267.905 118.025 268.105 118.755 ;
      RECT 268.4 118.025 268.6 118.755 ;
      RECT 269.22 118.025 269.42 118.755 ;
      RECT 269.715 118.025 269.915 118.755 ;
      RECT 270.215 118.025 270.415 118.755 ;
      RECT 270.37 0.52 270.63 2.335 ;
      RECT 270.715 118.025 270.915 118.755 ;
      RECT 270.88 0.52 271.14 14.11 ;
      RECT 271.21 118.025 271.41 118.755 ;
      RECT 272.255 0.17 273.025 0.94 ;
      RECT 272.765 0.17 273.025 8.7 ;
      RECT 272.255 0.17 272.515 12.9 ;
      RECT 271.745 0.52 272.005 2.485 ;
      RECT 272.03 118.025 272.23 118.755 ;
      RECT 273.275 0.17 274.045 0.43 ;
      RECT 273.785 0.17 274.045 10.48 ;
      RECT 273.275 0.17 273.535 10.99 ;
      RECT 272.525 118.025 272.725 118.755 ;
      RECT 273.025 118.025 273.225 118.755 ;
      RECT 273.525 118.025 273.725 118.755 ;
      RECT 274.02 118.025 274.22 118.755 ;
      RECT 275.315 0.17 276.085 0.43 ;
      RECT 275.315 0.17 275.575 11.5 ;
      RECT 275.825 0.17 276.085 11.5 ;
      RECT 274.84 118.025 275.04 118.755 ;
      RECT 275.335 118.025 275.535 118.755 ;
      RECT 276.335 0.17 277.105 0.94 ;
      RECT 276.335 0.17 276.595 12.9 ;
      RECT 276.845 0.17 277.105 12.9 ;
      RECT 275.835 118.025 276.035 118.755 ;
      RECT 276.335 118.025 276.535 118.755 ;
      RECT 276.83 118.025 277.03 118.755 ;
      RECT 277.355 0.52 277.615 5.815 ;
      RECT 278.21 0.52 278.47 5.16 ;
      RECT 278.21 4.9 278.99 5.16 ;
      RECT 278.73 4.9 278.99 6.64 ;
      RECT 277.65 118.025 277.85 118.755 ;
      RECT 278.145 118.025 278.345 118.755 ;
      RECT 278.645 118.025 278.845 118.755 ;
      RECT 279.145 118.025 279.345 118.755 ;
      RECT 279.64 118.025 279.84 118.755 ;
      RECT 280.46 118.025 280.66 118.755 ;
      RECT 280.955 118.025 281.155 118.755 ;
      RECT 281.455 118.025 281.655 118.755 ;
      RECT 281.61 0.52 281.87 2.335 ;
      RECT 281.955 118.025 282.155 118.755 ;
      RECT 282.12 0.52 282.38 14.11 ;
      RECT 282.45 118.025 282.65 118.755 ;
      RECT 283.495 0.17 284.265 0.94 ;
      RECT 284.005 0.17 284.265 8.7 ;
      RECT 283.495 0.17 283.755 12.9 ;
      RECT 282.985 0.52 283.245 2.485 ;
      RECT 283.27 118.025 283.47 118.755 ;
      RECT 284.515 0.17 285.285 0.43 ;
      RECT 285.025 0.17 285.285 10.48 ;
      RECT 284.515 0.17 284.775 10.99 ;
      RECT 283.765 118.025 283.965 118.755 ;
      RECT 284.265 118.025 284.465 118.755 ;
      RECT 284.765 118.025 284.965 118.755 ;
      RECT 285.26 118.025 285.46 118.755 ;
      RECT 286.555 0.17 287.325 0.43 ;
      RECT 286.555 0.17 286.815 11.5 ;
      RECT 287.065 0.17 287.325 11.5 ;
      RECT 286.08 118.025 286.28 118.755 ;
      RECT 286.575 118.025 286.775 118.755 ;
      RECT 287.575 0.17 288.345 0.94 ;
      RECT 287.575 0.17 287.835 12.9 ;
      RECT 288.085 0.17 288.345 12.9 ;
      RECT 287.075 118.025 287.275 118.755 ;
      RECT 287.575 118.025 287.775 118.755 ;
      RECT 288.07 118.025 288.27 118.755 ;
      RECT 288.595 0.52 288.855 5.815 ;
      RECT 289.45 0.52 289.71 5.16 ;
      RECT 289.45 4.9 290.23 5.16 ;
      RECT 289.97 4.9 290.23 6.64 ;
      RECT 288.89 118.025 289.09 118.755 ;
      RECT 289.385 118.025 289.585 118.755 ;
      RECT 289.885 118.025 290.085 118.755 ;
      RECT 290.385 118.025 290.585 118.755 ;
      RECT 290.88 118.025 291.08 118.755 ;
      RECT 291.7 118.025 291.9 118.755 ;
      RECT 292.195 118.025 292.395 118.755 ;
      RECT 292.695 118.025 292.895 118.755 ;
      RECT 292.85 0.52 293.11 2.335 ;
      RECT 293.195 118.025 293.395 118.755 ;
      RECT 293.36 0.52 293.62 14.11 ;
      RECT 293.69 118.025 293.89 118.755 ;
      RECT 294.735 0.17 295.505 0.94 ;
      RECT 295.245 0.17 295.505 8.7 ;
      RECT 294.735 0.17 294.995 12.9 ;
      RECT 294.225 0.52 294.485 2.485 ;
      RECT 294.51 118.025 294.71 118.755 ;
      RECT 295.755 0.17 296.525 0.43 ;
      RECT 296.265 0.17 296.525 10.48 ;
      RECT 295.755 0.17 296.015 10.99 ;
      RECT 295.005 118.025 295.205 118.755 ;
      RECT 295.505 118.025 295.705 118.755 ;
      RECT 296.005 118.025 296.205 118.755 ;
      RECT 296.5 118.025 296.7 118.755 ;
      RECT 297.795 0.17 298.565 0.43 ;
      RECT 297.795 0.17 298.055 11.5 ;
      RECT 298.305 0.17 298.565 11.5 ;
      RECT 297.32 118.025 297.52 118.755 ;
      RECT 297.815 118.025 298.015 118.755 ;
      RECT 298.815 0.17 299.585 0.94 ;
      RECT 298.815 0.17 299.075 12.9 ;
      RECT 299.325 0.17 299.585 12.9 ;
      RECT 298.315 118.025 298.515 118.755 ;
      RECT 298.815 118.025 299.015 118.755 ;
      RECT 299.31 118.025 299.51 118.755 ;
      RECT 299.835 0.52 300.095 5.815 ;
      RECT 300.69 0.52 300.95 5.16 ;
      RECT 300.69 4.9 301.47 5.16 ;
      RECT 301.21 4.9 301.47 6.64 ;
      RECT 300.13 118.025 300.33 118.755 ;
      RECT 300.625 118.025 300.825 118.755 ;
      RECT 301.125 118.025 301.325 118.755 ;
      RECT 301.625 118.025 301.825 118.755 ;
      RECT 302.12 118.025 302.32 118.755 ;
      RECT 302.94 118.025 303.14 118.755 ;
      RECT 303.435 118.025 303.635 118.755 ;
      RECT 303.935 118.025 304.135 118.755 ;
      RECT 304.09 0.52 304.35 2.335 ;
      RECT 304.435 118.025 304.635 118.755 ;
      RECT 304.6 0.52 304.86 14.11 ;
      RECT 304.93 118.025 305.13 118.755 ;
      RECT 305.975 0.17 306.745 0.94 ;
      RECT 306.485 0.17 306.745 8.7 ;
      RECT 305.975 0.17 306.235 12.9 ;
      RECT 305.465 0.52 305.725 2.485 ;
      RECT 305.75 118.025 305.95 118.755 ;
      RECT 306.995 0.17 307.765 0.43 ;
      RECT 307.505 0.17 307.765 10.48 ;
      RECT 306.995 0.17 307.255 10.99 ;
      RECT 306.245 118.025 306.445 118.755 ;
      RECT 306.745 118.025 306.945 118.755 ;
      RECT 307.245 118.025 307.445 118.755 ;
      RECT 307.74 118.025 307.94 118.755 ;
      RECT 309.035 0.17 309.805 0.43 ;
      RECT 309.035 0.17 309.295 11.5 ;
      RECT 309.545 0.17 309.805 11.5 ;
      RECT 308.56 118.025 308.76 118.755 ;
      RECT 309.055 118.025 309.255 118.755 ;
      RECT 310.055 0.17 310.825 0.94 ;
      RECT 310.055 0.17 310.315 12.9 ;
      RECT 310.565 0.17 310.825 12.9 ;
      RECT 309.555 118.025 309.755 118.755 ;
      RECT 310.055 118.025 310.255 118.755 ;
      RECT 310.55 118.025 310.75 118.755 ;
      RECT 311.075 0.52 311.335 5.815 ;
      RECT 311.93 0.52 312.19 5.16 ;
      RECT 311.93 4.9 312.71 5.16 ;
      RECT 312.45 4.9 312.71 6.64 ;
      RECT 311.37 118.025 311.57 118.755 ;
      RECT 311.865 118.025 312.065 118.755 ;
      RECT 312.365 118.025 312.565 118.755 ;
      RECT 312.865 118.025 313.065 118.755 ;
      RECT 313.36 118.025 313.56 118.755 ;
      RECT 314.18 118.025 314.38 118.755 ;
      RECT 314.675 118.025 314.875 118.755 ;
      RECT 315.175 118.025 315.375 118.755 ;
      RECT 315.33 0.52 315.59 2.335 ;
      RECT 315.675 118.025 315.875 118.755 ;
      RECT 315.84 0.52 316.1 14.11 ;
      RECT 316.17 118.025 316.37 118.755 ;
      RECT 317.215 0.17 317.985 0.94 ;
      RECT 317.725 0.17 317.985 8.7 ;
      RECT 317.215 0.17 317.475 12.9 ;
      RECT 316.705 0.52 316.965 2.485 ;
      RECT 316.99 118.025 317.19 118.755 ;
      RECT 318.235 0.17 319.005 0.43 ;
      RECT 318.745 0.17 319.005 10.48 ;
      RECT 318.235 0.17 318.495 10.99 ;
      RECT 317.485 118.025 317.685 118.755 ;
      RECT 317.985 118.025 318.185 118.755 ;
      RECT 318.485 118.025 318.685 118.755 ;
      RECT 318.98 118.025 319.18 118.755 ;
      RECT 320.275 0.17 321.045 0.43 ;
      RECT 320.275 0.17 320.535 11.5 ;
      RECT 320.785 0.17 321.045 11.5 ;
      RECT 319.8 118.025 320 118.755 ;
      RECT 320.295 118.025 320.495 118.755 ;
      RECT 321.295 0.17 322.065 0.94 ;
      RECT 321.295 0.17 321.555 12.9 ;
      RECT 321.805 0.17 322.065 12.9 ;
      RECT 320.795 118.025 320.995 118.755 ;
      RECT 321.295 118.025 321.495 118.755 ;
      RECT 321.79 118.025 321.99 118.755 ;
      RECT 322.315 0.52 322.575 5.815 ;
      RECT 323.17 0.52 323.43 5.16 ;
      RECT 323.17 4.9 323.95 5.16 ;
      RECT 323.69 4.9 323.95 6.64 ;
      RECT 322.61 118.025 322.81 118.755 ;
      RECT 323.105 118.025 323.305 118.755 ;
      RECT 323.605 118.025 323.805 118.755 ;
      RECT 324.105 118.025 324.305 118.755 ;
      RECT 324.6 118.025 324.8 118.755 ;
      RECT 325.42 118.025 325.62 118.755 ;
      RECT 325.915 118.025 326.115 118.755 ;
      RECT 326.415 118.025 326.615 118.755 ;
      RECT 326.57 0.52 326.83 2.335 ;
      RECT 326.915 118.025 327.115 118.755 ;
      RECT 327.08 0.52 327.34 14.11 ;
      RECT 327.41 118.025 327.61 118.755 ;
      RECT 328.455 0.17 329.225 0.94 ;
      RECT 328.965 0.17 329.225 8.7 ;
      RECT 328.455 0.17 328.715 12.9 ;
      RECT 327.945 0.52 328.205 2.485 ;
      RECT 328.23 118.025 328.43 118.755 ;
      RECT 329.475 0.17 330.245 0.43 ;
      RECT 329.985 0.17 330.245 10.48 ;
      RECT 329.475 0.17 329.735 10.99 ;
      RECT 328.725 118.025 328.925 118.755 ;
      RECT 329.225 118.025 329.425 118.755 ;
      RECT 329.725 118.025 329.925 118.755 ;
      RECT 330.22 118.025 330.42 118.755 ;
      RECT 331.515 0.17 332.285 0.43 ;
      RECT 331.515 0.17 331.775 11.5 ;
      RECT 332.025 0.17 332.285 11.5 ;
      RECT 331.04 118.025 331.24 118.755 ;
      RECT 331.535 118.025 331.735 118.755 ;
      RECT 332.535 0.17 333.305 0.94 ;
      RECT 332.535 0.17 332.795 12.9 ;
      RECT 333.045 0.17 333.305 12.9 ;
      RECT 332.035 118.025 332.235 118.755 ;
      RECT 332.535 118.025 332.735 118.755 ;
      RECT 333.03 118.025 333.23 118.755 ;
      RECT 333.555 0.52 333.815 5.815 ;
      RECT 334.41 0.52 334.67 5.16 ;
      RECT 334.41 4.9 335.19 5.16 ;
      RECT 334.93 4.9 335.19 6.64 ;
      RECT 333.85 118.025 334.05 118.755 ;
      RECT 334.345 118.025 334.545 118.755 ;
      RECT 334.845 118.025 335.045 118.755 ;
      RECT 335.345 118.025 335.545 118.755 ;
      RECT 335.84 118.025 336.04 118.755 ;
      RECT 336.66 118.025 336.86 118.755 ;
      RECT 337.155 118.025 337.355 118.755 ;
      RECT 337.655 118.025 337.855 118.755 ;
      RECT 337.81 0.52 338.07 2.335 ;
      RECT 338.155 118.025 338.355 118.755 ;
      RECT 338.32 0.52 338.58 14.11 ;
      RECT 338.65 118.025 338.85 118.755 ;
      RECT 339.695 0.17 340.465 0.94 ;
      RECT 340.205 0.17 340.465 8.7 ;
      RECT 339.695 0.17 339.955 12.9 ;
      RECT 339.185 0.52 339.445 2.485 ;
      RECT 339.47 118.025 339.67 118.755 ;
      RECT 340.715 0.17 341.485 0.43 ;
      RECT 341.225 0.17 341.485 10.48 ;
      RECT 340.715 0.17 340.975 10.99 ;
      RECT 339.965 118.025 340.165 118.755 ;
      RECT 340.465 118.025 340.665 118.755 ;
      RECT 340.965 118.025 341.165 118.755 ;
      RECT 341.46 118.025 341.66 118.755 ;
      RECT 342.755 0.17 343.525 0.43 ;
      RECT 342.755 0.17 343.015 11.5 ;
      RECT 343.265 0.17 343.525 11.5 ;
      RECT 342.28 118.025 342.48 118.755 ;
      RECT 342.775 118.025 342.975 118.755 ;
      RECT 343.775 0.17 344.545 0.94 ;
      RECT 343.775 0.17 344.035 12.9 ;
      RECT 344.285 0.17 344.545 12.9 ;
      RECT 343.275 118.025 343.475 118.755 ;
      RECT 343.775 118.025 343.975 118.755 ;
      RECT 344.27 118.025 344.47 118.755 ;
      RECT 344.795 0.52 345.055 5.815 ;
      RECT 345.65 0.52 345.91 5.16 ;
      RECT 345.65 4.9 346.43 5.16 ;
      RECT 346.17 4.9 346.43 6.64 ;
      RECT 345.09 118.025 345.29 118.755 ;
      RECT 345.585 118.025 345.785 118.755 ;
      RECT 346.085 118.025 346.285 118.755 ;
      RECT 346.585 118.025 346.785 118.755 ;
      RECT 347.08 118.025 347.28 118.755 ;
      RECT 347.9 118.025 348.1 118.755 ;
      RECT 348.395 118.025 348.595 118.755 ;
      RECT 348.895 118.025 349.095 118.755 ;
      RECT 349.05 0.52 349.31 2.335 ;
      RECT 349.395 118.025 349.595 118.755 ;
      RECT 349.56 0.52 349.82 14.11 ;
      RECT 349.89 118.025 350.09 118.755 ;
      RECT 350.935 0.17 351.705 0.94 ;
      RECT 351.445 0.17 351.705 8.7 ;
      RECT 350.935 0.17 351.195 12.9 ;
      RECT 350.425 0.52 350.685 2.485 ;
      RECT 350.71 118.025 350.91 118.755 ;
      RECT 351.955 0.17 352.725 0.43 ;
      RECT 352.465 0.17 352.725 10.48 ;
      RECT 351.955 0.17 352.215 10.99 ;
      RECT 351.205 118.025 351.405 118.755 ;
      RECT 351.705 118.025 351.905 118.755 ;
      RECT 352.205 118.025 352.405 118.755 ;
      RECT 352.7 118.025 352.9 118.755 ;
      RECT 353.995 0.17 354.765 0.43 ;
      RECT 353.995 0.17 354.255 11.5 ;
      RECT 354.505 0.17 354.765 11.5 ;
      RECT 353.52 118.025 353.72 118.755 ;
      RECT 354.015 118.025 354.215 118.755 ;
      RECT 355.015 0.17 355.785 0.94 ;
      RECT 355.015 0.17 355.275 12.9 ;
      RECT 355.525 0.17 355.785 12.9 ;
      RECT 354.515 118.025 354.715 118.755 ;
      RECT 355.015 118.025 355.215 118.755 ;
      RECT 355.51 118.025 355.71 118.755 ;
      RECT 356.035 0.52 356.295 5.815 ;
      RECT 356.89 0.52 357.15 5.16 ;
      RECT 356.89 4.9 357.67 5.16 ;
      RECT 357.41 4.9 357.67 6.64 ;
      RECT 356.33 118.025 356.53 118.755 ;
      RECT 356.825 118.025 357.025 118.755 ;
      RECT 357.325 118.025 357.525 118.755 ;
      RECT 357.825 118.025 358.025 118.755 ;
      RECT 358.32 118.025 358.52 118.755 ;
      RECT 359.14 118.025 359.34 118.755 ;
      RECT 359.635 118.025 359.835 118.755 ;
      RECT 360.135 118.025 360.335 118.755 ;
      RECT 360.29 0.52 360.55 2.335 ;
      RECT 360.635 118.025 360.835 118.755 ;
      RECT 360.8 0.52 361.06 14.11 ;
      RECT 361.13 118.025 361.33 118.755 ;
      RECT 362.175 0.17 362.945 0.94 ;
      RECT 362.685 0.17 362.945 8.7 ;
      RECT 362.175 0.17 362.435 12.9 ;
      RECT 361.665 0.52 361.925 2.485 ;
      RECT 361.95 118.025 362.15 118.755 ;
      RECT 363.195 0.17 363.965 0.43 ;
      RECT 363.705 0.17 363.965 10.48 ;
      RECT 363.195 0.17 363.455 10.99 ;
      RECT 362.445 118.025 362.645 118.755 ;
      RECT 362.945 118.025 363.145 118.755 ;
      RECT 363.445 118.025 363.645 118.755 ;
      RECT 363.94 118.025 364.14 118.755 ;
      RECT 365.235 0.17 366.005 0.43 ;
      RECT 365.235 0.17 365.495 11.5 ;
      RECT 365.745 0.17 366.005 11.5 ;
      RECT 364.76 118.025 364.96 118.755 ;
      RECT 365.255 118.025 365.455 118.755 ;
      RECT 366.255 0.17 367.025 0.94 ;
      RECT 366.255 0.17 366.515 12.9 ;
      RECT 366.765 0.17 367.025 12.9 ;
      RECT 365.755 118.025 365.955 118.755 ;
      RECT 366.255 118.025 366.455 118.755 ;
      RECT 366.75 118.025 366.95 118.755 ;
      RECT 367.275 0.52 367.535 5.815 ;
      RECT 368.13 0.52 368.39 5.16 ;
      RECT 368.13 4.9 368.91 5.16 ;
      RECT 368.65 4.9 368.91 6.64 ;
      RECT 367.57 118.025 367.77 118.755 ;
      RECT 368.065 118.025 368.265 118.755 ;
      RECT 368.565 118.025 368.765 118.755 ;
      RECT 369.065 118.025 369.265 118.755 ;
      RECT 369.56 118.025 369.76 118.755 ;
      RECT 370.38 118.025 370.58 118.755 ;
      RECT 370.875 118.025 371.075 118.755 ;
      RECT 371.375 118.025 371.575 118.755 ;
      RECT 371.53 0.52 371.79 2.335 ;
      RECT 371.875 118.025 372.075 118.755 ;
      RECT 372.04 0.52 372.3 14.11 ;
      RECT 372.37 118.025 372.57 118.755 ;
      RECT 373.415 0.17 374.185 0.94 ;
      RECT 373.925 0.17 374.185 8.7 ;
      RECT 373.415 0.17 373.675 12.9 ;
      RECT 372.905 0.52 373.165 2.485 ;
      RECT 373.19 118.025 373.39 118.755 ;
      RECT 374.435 0.17 375.205 0.43 ;
      RECT 374.945 0.17 375.205 10.48 ;
      RECT 374.435 0.17 374.695 10.99 ;
      RECT 373.685 118.025 373.885 118.755 ;
      RECT 374.185 118.025 374.385 118.755 ;
      RECT 374.685 118.025 374.885 118.755 ;
      RECT 375.18 118.025 375.38 118.755 ;
      RECT 376.475 0.17 377.245 0.43 ;
      RECT 376.475 0.17 376.735 11.5 ;
      RECT 376.985 0.17 377.245 11.5 ;
      RECT 376 118.025 376.2 118.755 ;
      RECT 376.495 118.025 376.695 118.755 ;
      RECT 377.495 0.17 378.265 0.94 ;
      RECT 377.495 0.17 377.755 12.9 ;
      RECT 378.005 0.17 378.265 12.9 ;
      RECT 376.995 118.025 377.195 118.755 ;
      RECT 377.495 118.025 377.695 118.755 ;
      RECT 377.99 118.025 378.19 118.755 ;
      RECT 378.515 0.52 378.775 5.815 ;
      RECT 379.37 0.52 379.63 5.16 ;
      RECT 379.37 4.9 380.15 5.16 ;
      RECT 379.89 4.9 380.15 6.64 ;
      RECT 378.81 118.025 379.01 118.755 ;
      RECT 379.305 118.025 379.505 118.755 ;
      RECT 379.805 118.025 380.005 118.755 ;
      RECT 380.305 118.025 380.505 118.755 ;
      RECT 380.8 118.025 381 118.755 ;
      RECT 381.62 118.025 381.82 118.755 ;
      RECT 382.115 118.025 382.315 118.755 ;
      RECT 382.615 118.025 382.815 118.755 ;
      RECT 382.77 0.52 383.03 2.335 ;
      RECT 383.115 118.025 383.315 118.755 ;
      RECT 383.28 0.52 383.54 14.11 ;
      RECT 383.61 118.025 383.81 118.755 ;
      RECT 384.655 0.17 385.425 0.94 ;
      RECT 385.165 0.17 385.425 8.7 ;
      RECT 384.655 0.17 384.915 12.9 ;
      RECT 384.145 0.52 384.405 2.485 ;
      RECT 384.43 118.025 384.63 118.755 ;
      RECT 385.675 0.17 386.445 0.43 ;
      RECT 386.185 0.17 386.445 10.48 ;
      RECT 385.675 0.17 385.935 10.99 ;
      RECT 384.925 118.025 385.125 118.755 ;
      RECT 385.425 118.025 385.625 118.755 ;
      RECT 385.925 118.025 386.125 118.755 ;
      RECT 386.42 118.025 386.62 118.755 ;
      RECT 387.715 0.17 388.485 0.43 ;
      RECT 387.715 0.17 387.975 11.5 ;
      RECT 388.225 0.17 388.485 11.5 ;
      RECT 387.24 118.025 387.44 118.755 ;
      RECT 387.735 118.025 387.935 118.755 ;
      RECT 388.735 0.17 389.505 0.94 ;
      RECT 388.735 0.17 388.995 12.9 ;
      RECT 389.245 0.17 389.505 12.9 ;
      RECT 388.235 118.025 388.435 118.755 ;
      RECT 388.735 118.025 388.935 118.755 ;
      RECT 389.23 118.025 389.43 118.755 ;
      RECT 389.755 0.52 390.015 5.815 ;
      RECT 390.61 0.52 390.87 5.16 ;
      RECT 390.61 4.9 391.39 5.16 ;
      RECT 391.13 4.9 391.39 6.64 ;
      RECT 390.05 118.025 390.25 118.755 ;
      RECT 390.545 118.025 390.745 118.755 ;
      RECT 391.045 118.025 391.245 118.755 ;
      RECT 391.545 118.025 391.745 118.755 ;
      RECT 392.04 118.025 392.24 118.755 ;
      RECT 392.86 118.025 393.06 118.755 ;
      RECT 393.355 118.025 393.555 118.755 ;
      RECT 393.855 118.025 394.055 118.755 ;
      RECT 394.01 0.52 394.27 2.335 ;
      RECT 394.355 118.025 394.555 118.755 ;
      RECT 394.52 0.52 394.78 14.11 ;
      RECT 394.85 118.025 395.05 118.755 ;
      RECT 395.895 0.17 396.665 0.94 ;
      RECT 396.405 0.17 396.665 8.7 ;
      RECT 395.895 0.17 396.155 12.9 ;
      RECT 395.385 0.52 395.645 2.485 ;
      RECT 395.67 118.025 395.87 118.755 ;
      RECT 396.915 0.17 397.685 0.43 ;
      RECT 397.425 0.17 397.685 10.48 ;
      RECT 396.915 0.17 397.175 10.99 ;
      RECT 396.165 118.025 396.365 118.755 ;
      RECT 396.665 118.025 396.865 118.755 ;
      RECT 397.165 118.025 397.365 118.755 ;
      RECT 397.66 118.025 397.86 118.755 ;
      RECT 398.955 0.17 399.725 0.43 ;
      RECT 398.955 0.17 399.215 11.5 ;
      RECT 399.465 0.17 399.725 11.5 ;
      RECT 398.48 118.025 398.68 118.755 ;
      RECT 398.975 118.025 399.175 118.755 ;
      RECT 399.975 0.17 400.745 0.94 ;
      RECT 399.975 0.17 400.235 12.9 ;
      RECT 400.485 0.17 400.745 12.9 ;
      RECT 399.475 118.025 399.675 118.755 ;
      RECT 399.975 118.025 400.175 118.755 ;
      RECT 400.47 118.025 400.67 118.755 ;
      RECT 400.995 0.52 401.255 5.815 ;
      RECT 401.85 0.52 402.11 5.16 ;
      RECT 401.85 4.9 402.63 5.16 ;
      RECT 402.37 4.9 402.63 6.64 ;
      RECT 401.29 118.025 401.49 118.755 ;
      RECT 401.785 118.025 401.985 118.755 ;
      RECT 402.285 118.025 402.485 118.755 ;
      RECT 402.785 118.025 402.985 118.755 ;
      RECT 403.28 118.025 403.48 118.755 ;
      RECT 404.1 118.025 404.3 118.755 ;
      RECT 404.595 118.025 404.795 118.755 ;
      RECT 405.095 118.025 405.295 118.755 ;
      RECT 405.25 0.52 405.51 2.335 ;
      RECT 405.595 118.025 405.795 118.755 ;
      RECT 405.76 0.52 406.02 14.11 ;
      RECT 406.09 118.025 406.29 118.755 ;
      RECT 407.135 0.17 407.905 0.94 ;
      RECT 407.645 0.17 407.905 8.7 ;
      RECT 407.135 0.17 407.395 12.9 ;
      RECT 406.625 0.52 406.885 2.485 ;
      RECT 406.91 118.025 407.11 118.755 ;
      RECT 408.155 0.17 408.925 0.43 ;
      RECT 408.665 0.17 408.925 10.48 ;
      RECT 408.155 0.17 408.415 10.99 ;
      RECT 407.405 118.025 407.605 118.755 ;
      RECT 407.905 118.025 408.105 118.755 ;
      RECT 408.405 118.025 408.605 118.755 ;
      RECT 408.9 118.025 409.1 118.755 ;
      RECT 410.195 0.17 410.965 0.43 ;
      RECT 410.195 0.17 410.455 11.5 ;
      RECT 410.705 0.17 410.965 11.5 ;
      RECT 409.72 118.025 409.92 118.755 ;
      RECT 410.215 118.025 410.415 118.755 ;
      RECT 411.215 0.17 411.985 0.94 ;
      RECT 411.215 0.17 411.475 12.9 ;
      RECT 411.725 0.17 411.985 12.9 ;
      RECT 410.715 118.025 410.915 118.755 ;
      RECT 411.215 118.025 411.415 118.755 ;
      RECT 411.71 118.025 411.91 118.755 ;
      RECT 412.235 0.52 412.495 5.815 ;
      RECT 413.09 0.52 413.35 5.16 ;
      RECT 413.09 4.9 413.87 5.16 ;
      RECT 413.61 4.9 413.87 6.64 ;
      RECT 412.53 118.025 412.73 118.755 ;
      RECT 413.025 118.025 413.225 118.755 ;
      RECT 413.525 118.025 413.725 118.755 ;
      RECT 414.025 118.025 414.225 118.755 ;
      RECT 414.52 118.025 414.72 118.755 ;
      RECT 415.34 118.025 415.54 118.755 ;
      RECT 416.335 45.465 416.535 118.755 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 194.32 0 200.69 118.78 ;
      RECT 209.63 0 210.89 118.78 ;
      RECT 238.545 0 243.375 118.78 ;
      RECT 249.785 0 254.615 118.78 ;
      RECT 261.025 0 265.855 118.78 ;
      RECT 272.265 0 277.095 118.78 ;
      RECT 283.505 0 288.335 118.78 ;
      RECT 294.745 0 299.575 118.78 ;
      RECT 305.985 0 310.815 118.78 ;
      RECT 317.225 0 322.055 118.78 ;
      RECT 328.465 0 333.295 118.78 ;
      RECT 339.705 0 344.535 118.78 ;
      RECT 350.945 0 355.775 118.78 ;
      RECT 362.185 0 367.015 118.78 ;
      RECT 373.425 0 378.255 118.78 ;
      RECT 384.665 0 389.495 118.78 ;
      RECT 395.905 0 400.735 118.78 ;
      RECT 407.145 0 411.975 118.78 ;
      RECT 201.98 0 202.22 118.78 ;
      RECT 203.51 0 203.75 118.78 ;
      RECT 206.57 0 206.81 118.78 ;
      RECT 208.1 0 208.34 118.78 ;
      RECT 215.23 0 224.15 118.78 ;
      RECT 0 0 3.03 118.78 ;
      RECT 4.655 0.17 9.505 118.78 ;
      RECT 11.65 0 14.27 118.78 ;
      RECT 15.895 0.17 20.745 118.78 ;
      RECT 22.89 0 25.51 118.78 ;
      RECT 27.135 0.17 31.985 118.78 ;
      RECT 34.13 0 36.75 118.78 ;
      RECT 38.375 0.17 43.225 118.78 ;
      RECT 45.37 0 47.99 118.78 ;
      RECT 49.615 0.17 54.465 118.78 ;
      RECT 56.61 0 59.23 118.78 ;
      RECT 60.855 0.17 65.705 118.78 ;
      RECT 67.85 0 70.47 118.78 ;
      RECT 72.095 0.17 76.945 118.78 ;
      RECT 79.09 0 81.71 118.78 ;
      RECT 83.335 0.17 88.185 118.78 ;
      RECT 90.33 0 92.95 118.78 ;
      RECT 94.575 0.17 99.425 118.78 ;
      RECT 101.57 0 104.19 118.78 ;
      RECT 105.815 0.17 110.665 118.78 ;
      RECT 112.81 0 115.43 118.78 ;
      RECT 117.055 0.17 121.905 118.78 ;
      RECT 124.05 0 126.67 118.78 ;
      RECT 128.295 0.17 133.145 118.78 ;
      RECT 135.29 0 137.91 118.78 ;
      RECT 139.535 0.17 144.385 118.78 ;
      RECT 146.53 0 149.15 118.78 ;
      RECT 150.775 0.17 155.625 118.78 ;
      RECT 157.77 0 160.39 118.78 ;
      RECT 162.015 0.17 166.865 118.78 ;
      RECT 169.01 0 171.63 118.78 ;
      RECT 173.255 0.17 178.105 118.78 ;
      RECT 180.25 0 192.03 118.78 ;
      RECT 194.32 0.17 200.7 118.78 ;
      RECT 201.97 0.3 202.23 118.78 ;
      RECT 203.5 0.3 203.76 118.78 ;
      RECT 206.56 0.3 206.82 118.78 ;
      RECT 208.09 0.3 208.35 118.78 ;
      RECT 209.63 0.17 210.9 118.78 ;
      RECT 209.62 0.3 210.9 118.78 ;
      RECT 215.23 0.3 224.16 118.78 ;
      RECT 224.93 0 236.39 118.78 ;
      RECT 224.92 0.17 236.39 118.78 ;
      RECT 238.535 0.17 243.385 118.78 ;
      RECT 245.01 0 247.63 118.78 ;
      RECT 249.775 0.17 254.625 118.78 ;
      RECT 256.25 0 258.87 118.78 ;
      RECT 261.015 0.17 265.865 118.78 ;
      RECT 267.49 0 270.11 118.78 ;
      RECT 272.255 0.17 277.105 118.78 ;
      RECT 278.73 0 281.35 118.78 ;
      RECT 283.495 0.17 288.345 118.78 ;
      RECT 289.97 0 292.59 118.78 ;
      RECT 294.735 0.17 299.585 118.78 ;
      RECT 301.21 0 303.83 118.78 ;
      RECT 305.975 0.17 310.825 118.78 ;
      RECT 312.45 0 315.07 118.78 ;
      RECT 317.215 0.17 322.065 118.78 ;
      RECT 323.69 0 326.31 118.78 ;
      RECT 328.455 0.17 333.305 118.78 ;
      RECT 334.93 0 337.55 118.78 ;
      RECT 339.695 0.17 344.545 118.78 ;
      RECT 346.17 0 348.79 118.78 ;
      RECT 350.935 0.17 355.785 118.78 ;
      RECT 357.41 0 360.03 118.78 ;
      RECT 362.175 0.17 367.025 118.78 ;
      RECT 368.65 0 371.27 118.78 ;
      RECT 373.415 0.17 378.265 118.78 ;
      RECT 379.89 0 382.51 118.78 ;
      RECT 384.655 0.17 389.505 118.78 ;
      RECT 391.13 0 393.75 118.78 ;
      RECT 395.895 0.17 400.745 118.78 ;
      RECT 402.37 0 404.99 118.78 ;
      RECT 407.135 0.17 411.985 118.78 ;
      RECT 413.61 0 416.64 118.78 ;
      RECT 0 0.52 416.64 118.78 ;
      RECT 4.665 0 9.495 118.78 ;
      RECT 15.905 0 20.735 118.78 ;
      RECT 27.145 0 31.975 118.78 ;
      RECT 38.385 0 43.215 118.78 ;
      RECT 49.625 0 54.455 118.78 ;
      RECT 60.865 0 65.695 118.78 ;
      RECT 72.105 0 76.935 118.78 ;
      RECT 83.345 0 88.175 118.78 ;
      RECT 94.585 0 99.415 118.78 ;
      RECT 105.825 0 110.655 118.78 ;
      RECT 117.065 0 121.895 118.78 ;
      RECT 128.305 0 133.135 118.78 ;
      RECT 139.545 0 144.375 118.78 ;
      RECT 150.785 0 155.615 118.78 ;
      RECT 162.025 0 166.855 118.78 ;
      RECT 173.265 0 178.095 118.78 ;
    LAYER Metal3 ;
      RECT 0 0 416.64 118.78 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 39.085 9.62 45.205 ;
      RECT 0 0 4 118.78 ;
      RECT 7.33 0 9.62 118.78 ;
      RECT 12.95 39.085 20.86 45.205 ;
      RECT 12.95 0 15.24 118.78 ;
      RECT 18.57 0 20.86 118.78 ;
      RECT 24.19 39.085 32.1 45.205 ;
      RECT 24.19 0 26.48 118.78 ;
      RECT 29.81 0 32.1 118.78 ;
      RECT 35.43 39.085 43.34 45.205 ;
      RECT 35.43 0 37.72 118.78 ;
      RECT 41.05 0 43.34 118.78 ;
      RECT 46.67 39.085 54.58 45.205 ;
      RECT 46.67 0 48.96 118.78 ;
      RECT 52.29 0 54.58 118.78 ;
      RECT 57.91 39.085 65.82 45.205 ;
      RECT 57.91 0 60.2 118.78 ;
      RECT 63.53 0 65.82 118.78 ;
      RECT 69.15 39.085 77.06 45.205 ;
      RECT 69.15 0 71.44 118.78 ;
      RECT 74.77 0 77.06 118.78 ;
      RECT 80.39 39.085 88.3 45.205 ;
      RECT 80.39 0 82.68 118.78 ;
      RECT 86.01 0 88.3 118.78 ;
      RECT 91.63 39.085 99.54 45.205 ;
      RECT 91.63 0 93.92 118.78 ;
      RECT 97.25 0 99.54 118.78 ;
      RECT 102.87 39.085 110.78 45.205 ;
      RECT 102.87 0 105.16 118.78 ;
      RECT 108.49 0 110.78 118.78 ;
      RECT 114.11 39.085 122.02 45.205 ;
      RECT 114.11 0 116.4 118.78 ;
      RECT 119.73 0 122.02 118.78 ;
      RECT 125.35 39.085 133.26 45.205 ;
      RECT 125.35 0 127.64 118.78 ;
      RECT 130.97 0 133.26 118.78 ;
      RECT 136.59 39.085 144.5 45.205 ;
      RECT 136.59 0 138.88 118.78 ;
      RECT 142.21 0 144.5 118.78 ;
      RECT 147.83 39.085 155.74 45.205 ;
      RECT 147.83 0 150.12 118.78 ;
      RECT 153.45 0 155.74 118.78 ;
      RECT 159.07 39.085 166.98 45.205 ;
      RECT 159.07 0 161.36 118.78 ;
      RECT 164.69 0 166.98 118.78 ;
      RECT 170.31 39.085 178.22 45.205 ;
      RECT 170.31 0 172.6 118.78 ;
      RECT 175.93 0 178.22 118.78 ;
      RECT 181.55 0 188.63 118.78 ;
      RECT 191.96 0 193.78 118.78 ;
      RECT 197.11 0 198.93 118.78 ;
      RECT 202.26 0 204.08 118.78 ;
      RECT 207.41 0 209.23 118.78 ;
      RECT 212.56 0 214.38 118.78 ;
      RECT 238.42 39.085 246.33 45.205 ;
      RECT 238.42 0 240.71 118.78 ;
      RECT 244.04 0 246.33 118.78 ;
      RECT 249.66 39.085 257.57 45.205 ;
      RECT 249.66 0 251.95 118.78 ;
      RECT 255.28 0 257.57 118.78 ;
      RECT 260.9 39.085 268.81 45.205 ;
      RECT 260.9 0 263.19 118.78 ;
      RECT 266.52 0 268.81 118.78 ;
      RECT 272.14 39.085 280.05 45.205 ;
      RECT 272.14 0 274.43 118.78 ;
      RECT 277.76 0 280.05 118.78 ;
      RECT 283.38 39.085 291.29 45.205 ;
      RECT 283.38 0 285.67 118.78 ;
      RECT 289 0 291.29 118.78 ;
      RECT 294.62 39.085 302.53 45.205 ;
      RECT 294.62 0 296.91 118.78 ;
      RECT 300.24 0 302.53 118.78 ;
      RECT 305.86 39.085 313.77 45.205 ;
      RECT 305.86 0 308.15 118.78 ;
      RECT 311.48 0 313.77 118.78 ;
      RECT 317.1 39.085 325.01 45.205 ;
      RECT 317.1 0 319.39 118.78 ;
      RECT 322.72 0 325.01 118.78 ;
      RECT 328.34 39.085 336.25 45.205 ;
      RECT 328.34 0 330.63 118.78 ;
      RECT 333.96 0 336.25 118.78 ;
      RECT 339.58 39.085 347.49 45.205 ;
      RECT 339.58 0 341.87 118.78 ;
      RECT 345.2 0 347.49 118.78 ;
      RECT 350.82 39.085 358.73 45.205 ;
      RECT 350.82 0 353.11 118.78 ;
      RECT 356.44 0 358.73 118.78 ;
      RECT 362.06 39.085 369.97 45.205 ;
      RECT 362.06 0 364.35 118.78 ;
      RECT 367.68 0 369.97 118.78 ;
      RECT 373.3 39.085 381.21 45.205 ;
      RECT 373.3 0 375.59 118.78 ;
      RECT 378.92 0 381.21 118.78 ;
      RECT 384.54 39.085 392.45 45.205 ;
      RECT 384.54 0 386.83 118.78 ;
      RECT 390.16 0 392.45 118.78 ;
      RECT 395.78 39.085 403.69 45.205 ;
      RECT 395.78 0 398.07 118.78 ;
      RECT 401.4 0 403.69 118.78 ;
      RECT 407.02 39.085 416.64 45.205 ;
      RECT 407.02 0 409.31 118.78 ;
      RECT 412.64 0 416.64 118.78 ;
      RECT 217.71 0 219.53 118.78 ;
      RECT 222.86 0 224.68 118.78 ;
      RECT 228.01 0 235.09 118.78 ;
  END
END RM_IHPSG13_1P_256x32_c2_bm_bist

END LIBRARY
