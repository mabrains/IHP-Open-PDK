# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 16:20:24 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_512x8_c3_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_512x8_c3_bm_bist 0 0 ;
  SIZE 236.8 BY 110.38 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.09 0 155.35 0.26 ;
    END
  END A_DIN[4]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.45 0 81.71 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.56 0 153.82 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.98 0 83.24 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.97 0 159.23 0.26 ;
    END
  END A_BM[4]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.57 0 77.83 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.5 0 160.76 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.04 0 76.3 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 159.835 0 160.095 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.705 0 76.965 0.26 ;
    END
  END A_DOUT[3]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 224.11 0 226.92 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.87 0 215.68 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 201.63 0 204.44 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.39 0 193.2 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.15 0 181.96 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.91 0 170.72 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.67 0 159.48 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.43 0 148.24 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.02 0 137.83 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.72 0 127.53 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.27 0 112.08 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 98.97 0 101.78 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 110.38 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 0 232.54 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 0 221.3 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 0 210.06 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 0 198.82 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 0 187.58 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 0 176.34 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 0 165.1 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 0 153.86 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.87 0 132.68 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.57 0 122.38 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.42 0 117.23 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 104.12 0 106.93 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 30.425 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 37.065 232.54 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 37.065 221.3 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 37.065 210.06 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 37.065 198.82 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 37.065 187.58 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 37.065 176.34 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 37.065 165.1 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 37.065 153.86 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 37.065 85.75 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 37.065 74.51 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 37.065 63.27 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 37.065 52.03 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 37.065 40.79 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 37.065 29.55 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 37.065 18.31 110.38 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 37.065 7.07 110.38 ;
    END
  END VDDARRAY!
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 177.57 0 177.83 0.26 ;
    END
  END A_DIN[5]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 58.97 0 59.23 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.04 0 176.3 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.5 0 60.76 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.45 0 181.71 0.26 ;
    END
  END A_BM[5]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.09 0 55.35 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.98 0 183.24 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.56 0 53.82 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.315 0 182.575 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.225 0 54.485 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.05 0 200.31 0.26 ;
    END
  END A_DIN[6]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.49 0 36.75 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 198.52 0 198.78 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.02 0 38.28 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.93 0 204.19 0.26 ;
    END
  END A_BM[6]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.61 0 32.87 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.46 0 205.72 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.08 0 31.34 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.795 0 205.055 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.745 0 32.005 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 222.53 0 222.79 0.26 ;
    END
  END A_DIN[7]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.01 0 14.27 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221 0 221.26 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.54 0 15.8 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.41 0 226.67 0.26 ;
    END
  END A_BM[7]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.13 0 10.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.94 0 228.2 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 8.6 0 8.86 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.275 0 227.535 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.265 0 9.525 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7171 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 34.349515 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.6 0 114.86 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5127 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 38.31068 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.19 0 119.45 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.59 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 28.783172 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.09 0 114.35 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3856 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 32.744337 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 118.68 0 118.94 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4519 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 33.029126 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.81 0 100.07 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1867 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 31.708738 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.34 0 101.6 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.25 0 122.51 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.76 0 123.02 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.23 0 121.49 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.74 0 122 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0139 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.763754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.8 0 125.06 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7487 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.443366 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.29 0 124.55 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7429 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 59.372168 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.78 0 124.04 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4777 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 58.05178 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.27 0 123.53 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.36 0 102.62 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4931 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.191934 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.87 0 103.13 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2323 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 51.851133 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.38 0 103.64 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9671 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.530744 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.89 0 104.15 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8707 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.220065 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.56 0 112.82 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81105 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.923077 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.13 0 116.39 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.62 0 115.88 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8407 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.09186 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.07 0 113.33 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.874 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 12.046332 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.49 0 134.75 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 72.69295 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.3675 LAYER Metal3 ;
      ANTENNAMAXAREACAR 1.686364 LAYER Metal2 ;
      ANTENNAMAXAREACAR 13.950709 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.11 0 115.37 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9799 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 11.079661 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.03 0 111.29 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9279 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.820762 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.66 0 117.92 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7211 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.812298 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.15 0 117.41 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7137 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.775454 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.54 0 111.8 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 236.8 110.38 ;
    LAYER Metal2 ;
      RECT 0.105 37.065 0.305 110.355 ;
      RECT 1.1 109.625 1.3 110.355 ;
      RECT 1.92 109.625 2.12 110.355 ;
      RECT 2.415 109.625 2.615 110.355 ;
      RECT 2.915 109.625 3.115 110.355 ;
      RECT 3.415 109.625 3.615 110.355 ;
      RECT 3.91 109.625 4.11 110.355 ;
      RECT 4.73 109.625 4.93 110.355 ;
      RECT 5.225 109.625 5.425 110.355 ;
      RECT 5.725 109.625 5.925 110.355 ;
      RECT 7.225 0.17 7.995 0.43 ;
      RECT 7.225 0.17 7.485 11.38 ;
      RECT 7.735 0.17 7.995 17.1 ;
      RECT 6.225 109.625 6.425 110.355 ;
      RECT 6.72 109.625 6.92 110.355 ;
      RECT 7.54 109.625 7.74 110.355 ;
      RECT 8.035 109.625 8.235 110.355 ;
      RECT 8.535 109.625 8.735 110.355 ;
      RECT 8.6 0.52 8.86 2.255 ;
      RECT 9.035 109.625 9.235 110.355 ;
      RECT 9.265 0.52 9.525 8.085 ;
      RECT 9.53 109.625 9.73 110.355 ;
      RECT 10.13 0.52 10.39 1.5 ;
      RECT 10.35 109.625 10.55 110.355 ;
      RECT 10.845 109.625 11.045 110.355 ;
      RECT 11.345 109.625 11.545 110.355 ;
      RECT 11.845 109.625 12.045 110.355 ;
      RECT 12.34 109.625 12.54 110.355 ;
      RECT 13.16 109.625 13.36 110.355 ;
      RECT 13.655 109.625 13.855 110.355 ;
      RECT 14.01 0.52 14.27 2.255 ;
      RECT 14.155 109.625 14.355 110.355 ;
      RECT 14.655 109.625 14.855 110.355 ;
      RECT 15.15 109.625 15.35 110.355 ;
      RECT 16.255 0.8 17.025 1.57 ;
      RECT 16.255 0.3 16.515 13.03 ;
      RECT 16.765 0.3 17.025 13.03 ;
      RECT 15.54 0.52 15.8 2.255 ;
      RECT 15.97 109.625 16.17 110.355 ;
      RECT 16.465 109.625 16.665 110.355 ;
      RECT 16.965 109.625 17.165 110.355 ;
      RECT 17.465 109.625 17.665 110.355 ;
      RECT 17.96 109.625 18.16 110.355 ;
      RECT 18.78 109.625 18.98 110.355 ;
      RECT 19.975 0.17 20.745 0.43 ;
      RECT 19.975 0.17 20.235 13.055 ;
      RECT 20.485 0.17 20.745 13.055 ;
      RECT 19.275 109.625 19.475 110.355 ;
      RECT 19.775 109.625 19.975 110.355 ;
      RECT 20.275 109.625 20.475 110.355 ;
      RECT 20.77 109.625 20.97 110.355 ;
      RECT 21.59 109.625 21.79 110.355 ;
      RECT 22.085 109.625 22.285 110.355 ;
      RECT 22.585 109.625 22.785 110.355 ;
      RECT 23.085 109.625 23.285 110.355 ;
      RECT 23.58 109.625 23.78 110.355 ;
      RECT 24.4 109.625 24.6 110.355 ;
      RECT 24.895 109.625 25.095 110.355 ;
      RECT 25.395 109.625 25.595 110.355 ;
      RECT 25.895 109.625 26.095 110.355 ;
      RECT 26.39 109.625 26.59 110.355 ;
      RECT 27.21 109.625 27.41 110.355 ;
      RECT 27.705 109.625 27.905 110.355 ;
      RECT 28.205 109.625 28.405 110.355 ;
      RECT 29.705 0.17 30.475 0.43 ;
      RECT 29.705 0.17 29.965 11.38 ;
      RECT 30.215 0.17 30.475 17.1 ;
      RECT 28.705 109.625 28.905 110.355 ;
      RECT 29.2 109.625 29.4 110.355 ;
      RECT 30.02 109.625 30.22 110.355 ;
      RECT 30.515 109.625 30.715 110.355 ;
      RECT 31.015 109.625 31.215 110.355 ;
      RECT 31.08 0.52 31.34 2.255 ;
      RECT 31.515 109.625 31.715 110.355 ;
      RECT 31.745 0.52 32.005 8.085 ;
      RECT 32.01 109.625 32.21 110.355 ;
      RECT 32.61 0.52 32.87 1.5 ;
      RECT 32.83 109.625 33.03 110.355 ;
      RECT 33.325 109.625 33.525 110.355 ;
      RECT 33.825 109.625 34.025 110.355 ;
      RECT 34.325 109.625 34.525 110.355 ;
      RECT 34.82 109.625 35.02 110.355 ;
      RECT 35.64 109.625 35.84 110.355 ;
      RECT 36.135 109.625 36.335 110.355 ;
      RECT 36.49 0.52 36.75 2.255 ;
      RECT 36.635 109.625 36.835 110.355 ;
      RECT 37.135 109.625 37.335 110.355 ;
      RECT 37.63 109.625 37.83 110.355 ;
      RECT 38.735 0.8 39.505 1.57 ;
      RECT 38.735 0.3 38.995 13.03 ;
      RECT 39.245 0.3 39.505 13.03 ;
      RECT 38.02 0.52 38.28 2.255 ;
      RECT 38.45 109.625 38.65 110.355 ;
      RECT 38.945 109.625 39.145 110.355 ;
      RECT 39.445 109.625 39.645 110.355 ;
      RECT 39.945 109.625 40.145 110.355 ;
      RECT 40.44 109.625 40.64 110.355 ;
      RECT 41.26 109.625 41.46 110.355 ;
      RECT 42.455 0.17 43.225 0.43 ;
      RECT 42.455 0.17 42.715 13.055 ;
      RECT 42.965 0.17 43.225 13.055 ;
      RECT 41.755 109.625 41.955 110.355 ;
      RECT 42.255 109.625 42.455 110.355 ;
      RECT 42.755 109.625 42.955 110.355 ;
      RECT 43.25 109.625 43.45 110.355 ;
      RECT 44.07 109.625 44.27 110.355 ;
      RECT 44.565 109.625 44.765 110.355 ;
      RECT 45.065 109.625 45.265 110.355 ;
      RECT 45.565 109.625 45.765 110.355 ;
      RECT 46.06 109.625 46.26 110.355 ;
      RECT 46.88 109.625 47.08 110.355 ;
      RECT 47.375 109.625 47.575 110.355 ;
      RECT 47.875 109.625 48.075 110.355 ;
      RECT 48.375 109.625 48.575 110.355 ;
      RECT 48.87 109.625 49.07 110.355 ;
      RECT 49.69 109.625 49.89 110.355 ;
      RECT 50.185 109.625 50.385 110.355 ;
      RECT 50.685 109.625 50.885 110.355 ;
      RECT 52.185 0.17 52.955 0.43 ;
      RECT 52.185 0.17 52.445 11.38 ;
      RECT 52.695 0.17 52.955 17.1 ;
      RECT 51.185 109.625 51.385 110.355 ;
      RECT 51.68 109.625 51.88 110.355 ;
      RECT 52.5 109.625 52.7 110.355 ;
      RECT 52.995 109.625 53.195 110.355 ;
      RECT 53.495 109.625 53.695 110.355 ;
      RECT 53.56 0.52 53.82 2.255 ;
      RECT 53.995 109.625 54.195 110.355 ;
      RECT 54.225 0.52 54.485 8.085 ;
      RECT 54.49 109.625 54.69 110.355 ;
      RECT 55.09 0.52 55.35 1.5 ;
      RECT 55.31 109.625 55.51 110.355 ;
      RECT 55.805 109.625 56.005 110.355 ;
      RECT 56.305 109.625 56.505 110.355 ;
      RECT 56.805 109.625 57.005 110.355 ;
      RECT 57.3 109.625 57.5 110.355 ;
      RECT 58.12 109.625 58.32 110.355 ;
      RECT 58.615 109.625 58.815 110.355 ;
      RECT 58.97 0.52 59.23 2.255 ;
      RECT 59.115 109.625 59.315 110.355 ;
      RECT 59.615 109.625 59.815 110.355 ;
      RECT 60.11 109.625 60.31 110.355 ;
      RECT 61.215 0.8 61.985 1.57 ;
      RECT 61.215 0.3 61.475 13.03 ;
      RECT 61.725 0.3 61.985 13.03 ;
      RECT 60.5 0.52 60.76 2.255 ;
      RECT 60.93 109.625 61.13 110.355 ;
      RECT 61.425 109.625 61.625 110.355 ;
      RECT 61.925 109.625 62.125 110.355 ;
      RECT 62.425 109.625 62.625 110.355 ;
      RECT 62.92 109.625 63.12 110.355 ;
      RECT 63.74 109.625 63.94 110.355 ;
      RECT 64.935 0.17 65.705 0.43 ;
      RECT 64.935 0.17 65.195 13.055 ;
      RECT 65.445 0.17 65.705 13.055 ;
      RECT 64.235 109.625 64.435 110.355 ;
      RECT 64.735 109.625 64.935 110.355 ;
      RECT 65.235 109.625 65.435 110.355 ;
      RECT 65.73 109.625 65.93 110.355 ;
      RECT 66.55 109.625 66.75 110.355 ;
      RECT 67.045 109.625 67.245 110.355 ;
      RECT 67.545 109.625 67.745 110.355 ;
      RECT 68.045 109.625 68.245 110.355 ;
      RECT 68.54 109.625 68.74 110.355 ;
      RECT 69.36 109.625 69.56 110.355 ;
      RECT 69.855 109.625 70.055 110.355 ;
      RECT 70.355 109.625 70.555 110.355 ;
      RECT 70.855 109.625 71.055 110.355 ;
      RECT 71.35 109.625 71.55 110.355 ;
      RECT 72.17 109.625 72.37 110.355 ;
      RECT 72.665 109.625 72.865 110.355 ;
      RECT 73.165 109.625 73.365 110.355 ;
      RECT 74.665 0.17 75.435 0.43 ;
      RECT 74.665 0.17 74.925 11.38 ;
      RECT 75.175 0.17 75.435 17.1 ;
      RECT 73.665 109.625 73.865 110.355 ;
      RECT 74.16 109.625 74.36 110.355 ;
      RECT 74.98 109.625 75.18 110.355 ;
      RECT 75.475 109.625 75.675 110.355 ;
      RECT 75.975 109.625 76.175 110.355 ;
      RECT 76.04 0.52 76.3 2.255 ;
      RECT 76.475 109.625 76.675 110.355 ;
      RECT 76.705 0.52 76.965 8.085 ;
      RECT 76.97 109.625 77.17 110.355 ;
      RECT 77.57 0.52 77.83 1.5 ;
      RECT 77.79 109.625 77.99 110.355 ;
      RECT 78.285 109.625 78.485 110.355 ;
      RECT 78.785 109.625 78.985 110.355 ;
      RECT 79.285 109.625 79.485 110.355 ;
      RECT 79.78 109.625 79.98 110.355 ;
      RECT 80.6 109.625 80.8 110.355 ;
      RECT 81.095 109.625 81.295 110.355 ;
      RECT 81.45 0.52 81.71 2.255 ;
      RECT 81.595 109.625 81.795 110.355 ;
      RECT 82.095 109.625 82.295 110.355 ;
      RECT 82.59 109.625 82.79 110.355 ;
      RECT 83.695 0.8 84.465 1.57 ;
      RECT 83.695 0.3 83.955 13.03 ;
      RECT 84.205 0.3 84.465 13.03 ;
      RECT 82.98 0.52 83.24 2.255 ;
      RECT 83.41 109.625 83.61 110.355 ;
      RECT 83.905 109.625 84.105 110.355 ;
      RECT 84.405 109.625 84.605 110.355 ;
      RECT 84.905 109.625 85.105 110.355 ;
      RECT 85.4 109.625 85.6 110.355 ;
      RECT 86.22 109.625 86.42 110.355 ;
      RECT 87.415 0.17 88.185 0.43 ;
      RECT 87.415 0.17 87.675 13.055 ;
      RECT 87.925 0.17 88.185 13.055 ;
      RECT 86.715 109.625 86.915 110.355 ;
      RECT 87.215 109.625 87.415 110.355 ;
      RECT 87.715 109.625 87.915 110.355 ;
      RECT 88.21 109.625 88.41 110.355 ;
      RECT 89.03 109.625 89.23 110.355 ;
      RECT 89.525 109.625 89.725 110.355 ;
      RECT 90.025 109.625 90.225 110.355 ;
      RECT 90.525 109.625 90.725 110.355 ;
      RECT 96.595 0.17 97.365 0.43 ;
      RECT 96.595 0.17 96.855 36.945 ;
      RECT 97.105 0.17 97.365 36.945 ;
      RECT 91.02 109.625 91.22 110.355 ;
      RECT 91.84 109.625 92.04 110.355 ;
      RECT 99.3 0 99.56 4.94 ;
      RECT 99.3 4.68 100.07 4.94 ;
      RECT 99.81 4.68 100.07 12.9 ;
      RECT 99.81 0.52 100.07 1.78 ;
      RECT 99.81 1.52 100.58 1.78 ;
      RECT 100.32 1.52 100.58 12.9 ;
      RECT 92.835 109.625 93.035 110.355 ;
      RECT 100.32 0.59 101.09 1.27 ;
      RECT 100.83 0.59 101.09 7.965 ;
      RECT 97.615 0.3 97.875 37.365 ;
      RECT 98.125 0.3 98.385 37.365 ;
      RECT 101.34 0.52 101.6 12.9 ;
      RECT 101.85 0 102.11 12.9 ;
      RECT 102.36 0.52 102.62 12.9 ;
      RECT 102.87 0.52 103.13 12.9 ;
      RECT 103.38 0.52 103.64 12.9 ;
      RECT 106.44 0.17 107.21 0.43 ;
      RECT 106.44 0.17 106.7 2.085 ;
      RECT 106.95 0.17 107.21 9 ;
      RECT 103.89 0.52 104.15 12.9 ;
      RECT 104.4 0 104.66 8.565 ;
      RECT 104.91 0 105.17 8.055 ;
      RECT 111.03 0.52 111.29 6.59 ;
      RECT 112.56 0.52 112.82 6.305 ;
      RECT 112.56 6.045 113.53 6.305 ;
      RECT 111.54 0.52 111.8 2.23 ;
      RECT 113.07 0.52 113.33 2.955 ;
      RECT 114.09 0.52 114.35 12.9 ;
      RECT 114.6 0.52 114.86 12.9 ;
      RECT 116.13 0.52 116.39 6.29 ;
      RECT 115.62 6.045 116.39 6.29 ;
      RECT 115.11 0.52 115.37 6.745 ;
      RECT 117.66 0.52 117.92 6.59 ;
      RECT 117.015 6.33 117.92 6.59 ;
      RECT 115.62 0.52 115.88 2.955 ;
      RECT 117.15 0.52 117.41 2.67 ;
      RECT 118.68 0.52 118.94 12.9 ;
      RECT 119.19 0.52 119.45 12.9 ;
      RECT 120.72 0.575 120.98 7.965 ;
      RECT 121.23 0.52 121.49 12.9 ;
      RECT 121.74 0.52 122 12.9 ;
      RECT 122.25 0.52 122.51 12.9 ;
      RECT 122.76 0.52 123.02 12.9 ;
      RECT 123.27 0.52 123.53 12.9 ;
      RECT 123.78 0.52 124.04 12.9 ;
      RECT 124.29 0.52 124.55 12.9 ;
      RECT 124.8 0.52 125.06 12.9 ;
      RECT 125.31 0 125.57 12.9 ;
      RECT 125.82 0 126.08 12.9 ;
      RECT 127.35 0 127.61 12.9 ;
      RECT 127.86 0 128.12 12.9 ;
      RECT 135 0.17 135.77 0.43 ;
      RECT 135 0.17 135.26 13.845 ;
      RECT 135.51 0.17 135.77 13.845 ;
      RECT 137.04 0.17 137.81 0.43 ;
      RECT 137.04 0.17 137.3 2.11 ;
      RECT 137.55 0.17 137.81 2.11 ;
      RECT 132.45 0 132.71 3.61 ;
      RECT 132.96 0 133.22 4.12 ;
      RECT 139.435 0.17 140.205 0.43 ;
      RECT 139.435 0.17 139.695 36.945 ;
      RECT 139.945 0.17 140.205 36.945 ;
      RECT 134.49 0.52 134.75 15.16 ;
      RECT 138.415 0.3 138.675 37.365 ;
      RECT 138.925 0.3 139.185 37.365 ;
      RECT 143.765 109.625 143.965 110.355 ;
      RECT 144.76 109.625 144.96 110.355 ;
      RECT 145.58 109.625 145.78 110.355 ;
      RECT 146.075 109.625 146.275 110.355 ;
      RECT 146.575 109.625 146.775 110.355 ;
      RECT 147.075 109.625 147.275 110.355 ;
      RECT 148.615 0.17 149.385 0.43 ;
      RECT 148.615 0.17 148.875 13.055 ;
      RECT 149.125 0.17 149.385 13.055 ;
      RECT 147.57 109.625 147.77 110.355 ;
      RECT 148.39 109.625 148.59 110.355 ;
      RECT 148.885 109.625 149.085 110.355 ;
      RECT 149.385 109.625 149.585 110.355 ;
      RECT 149.885 109.625 150.085 110.355 ;
      RECT 150.38 109.625 150.58 110.355 ;
      RECT 151.2 109.625 151.4 110.355 ;
      RECT 152.335 0.8 153.105 1.57 ;
      RECT 152.335 0.3 152.595 13.03 ;
      RECT 152.845 0.3 153.105 13.03 ;
      RECT 151.695 109.625 151.895 110.355 ;
      RECT 152.195 109.625 152.395 110.355 ;
      RECT 152.695 109.625 152.895 110.355 ;
      RECT 153.19 109.625 153.39 110.355 ;
      RECT 153.56 0.52 153.82 2.255 ;
      RECT 154.01 109.625 154.21 110.355 ;
      RECT 154.505 109.625 154.705 110.355 ;
      RECT 155.005 109.625 155.205 110.355 ;
      RECT 155.09 0.52 155.35 2.255 ;
      RECT 155.505 109.625 155.705 110.355 ;
      RECT 156 109.625 156.2 110.355 ;
      RECT 156.82 109.625 157.02 110.355 ;
      RECT 157.315 109.625 157.515 110.355 ;
      RECT 157.815 109.625 158.015 110.355 ;
      RECT 158.315 109.625 158.515 110.355 ;
      RECT 158.81 109.625 159.01 110.355 ;
      RECT 158.97 0.52 159.23 1.5 ;
      RECT 159.63 109.625 159.83 110.355 ;
      RECT 159.835 0.52 160.095 8.085 ;
      RECT 160.125 109.625 160.325 110.355 ;
      RECT 160.5 0.52 160.76 2.255 ;
      RECT 161.365 0.17 162.135 0.43 ;
      RECT 161.875 0.17 162.135 11.38 ;
      RECT 161.365 0.17 161.625 17.1 ;
      RECT 160.625 109.625 160.825 110.355 ;
      RECT 161.125 109.625 161.325 110.355 ;
      RECT 161.62 109.625 161.82 110.355 ;
      RECT 162.44 109.625 162.64 110.355 ;
      RECT 162.935 109.625 163.135 110.355 ;
      RECT 163.435 109.625 163.635 110.355 ;
      RECT 163.935 109.625 164.135 110.355 ;
      RECT 164.43 109.625 164.63 110.355 ;
      RECT 165.25 109.625 165.45 110.355 ;
      RECT 165.745 109.625 165.945 110.355 ;
      RECT 166.245 109.625 166.445 110.355 ;
      RECT 166.745 109.625 166.945 110.355 ;
      RECT 167.24 109.625 167.44 110.355 ;
      RECT 168.06 109.625 168.26 110.355 ;
      RECT 168.555 109.625 168.755 110.355 ;
      RECT 169.055 109.625 169.255 110.355 ;
      RECT 169.555 109.625 169.755 110.355 ;
      RECT 171.095 0.17 171.865 0.43 ;
      RECT 171.095 0.17 171.355 13.055 ;
      RECT 171.605 0.17 171.865 13.055 ;
      RECT 170.05 109.625 170.25 110.355 ;
      RECT 170.87 109.625 171.07 110.355 ;
      RECT 171.365 109.625 171.565 110.355 ;
      RECT 171.865 109.625 172.065 110.355 ;
      RECT 172.365 109.625 172.565 110.355 ;
      RECT 172.86 109.625 173.06 110.355 ;
      RECT 173.68 109.625 173.88 110.355 ;
      RECT 174.815 0.8 175.585 1.57 ;
      RECT 174.815 0.3 175.075 13.03 ;
      RECT 175.325 0.3 175.585 13.03 ;
      RECT 174.175 109.625 174.375 110.355 ;
      RECT 174.675 109.625 174.875 110.355 ;
      RECT 175.175 109.625 175.375 110.355 ;
      RECT 175.67 109.625 175.87 110.355 ;
      RECT 176.04 0.52 176.3 2.255 ;
      RECT 176.49 109.625 176.69 110.355 ;
      RECT 176.985 109.625 177.185 110.355 ;
      RECT 177.485 109.625 177.685 110.355 ;
      RECT 177.57 0.52 177.83 2.255 ;
      RECT 177.985 109.625 178.185 110.355 ;
      RECT 178.48 109.625 178.68 110.355 ;
      RECT 179.3 109.625 179.5 110.355 ;
      RECT 179.795 109.625 179.995 110.355 ;
      RECT 180.295 109.625 180.495 110.355 ;
      RECT 180.795 109.625 180.995 110.355 ;
      RECT 181.29 109.625 181.49 110.355 ;
      RECT 181.45 0.52 181.71 1.5 ;
      RECT 182.11 109.625 182.31 110.355 ;
      RECT 182.315 0.52 182.575 8.085 ;
      RECT 182.605 109.625 182.805 110.355 ;
      RECT 182.98 0.52 183.24 2.255 ;
      RECT 183.845 0.17 184.615 0.43 ;
      RECT 184.355 0.17 184.615 11.38 ;
      RECT 183.845 0.17 184.105 17.1 ;
      RECT 183.105 109.625 183.305 110.355 ;
      RECT 183.605 109.625 183.805 110.355 ;
      RECT 184.1 109.625 184.3 110.355 ;
      RECT 184.92 109.625 185.12 110.355 ;
      RECT 185.415 109.625 185.615 110.355 ;
      RECT 185.915 109.625 186.115 110.355 ;
      RECT 186.415 109.625 186.615 110.355 ;
      RECT 186.91 109.625 187.11 110.355 ;
      RECT 187.73 109.625 187.93 110.355 ;
      RECT 188.225 109.625 188.425 110.355 ;
      RECT 188.725 109.625 188.925 110.355 ;
      RECT 189.225 109.625 189.425 110.355 ;
      RECT 189.72 109.625 189.92 110.355 ;
      RECT 190.54 109.625 190.74 110.355 ;
      RECT 191.035 109.625 191.235 110.355 ;
      RECT 191.535 109.625 191.735 110.355 ;
      RECT 192.035 109.625 192.235 110.355 ;
      RECT 193.575 0.17 194.345 0.43 ;
      RECT 193.575 0.17 193.835 13.055 ;
      RECT 194.085 0.17 194.345 13.055 ;
      RECT 192.53 109.625 192.73 110.355 ;
      RECT 193.35 109.625 193.55 110.355 ;
      RECT 193.845 109.625 194.045 110.355 ;
      RECT 194.345 109.625 194.545 110.355 ;
      RECT 194.845 109.625 195.045 110.355 ;
      RECT 195.34 109.625 195.54 110.355 ;
      RECT 196.16 109.625 196.36 110.355 ;
      RECT 197.295 0.8 198.065 1.57 ;
      RECT 197.295 0.3 197.555 13.03 ;
      RECT 197.805 0.3 198.065 13.03 ;
      RECT 196.655 109.625 196.855 110.355 ;
      RECT 197.155 109.625 197.355 110.355 ;
      RECT 197.655 109.625 197.855 110.355 ;
      RECT 198.15 109.625 198.35 110.355 ;
      RECT 198.52 0.52 198.78 2.255 ;
      RECT 198.97 109.625 199.17 110.355 ;
      RECT 199.465 109.625 199.665 110.355 ;
      RECT 199.965 109.625 200.165 110.355 ;
      RECT 200.05 0.52 200.31 2.255 ;
      RECT 200.465 109.625 200.665 110.355 ;
      RECT 200.96 109.625 201.16 110.355 ;
      RECT 201.78 109.625 201.98 110.355 ;
      RECT 202.275 109.625 202.475 110.355 ;
      RECT 202.775 109.625 202.975 110.355 ;
      RECT 203.275 109.625 203.475 110.355 ;
      RECT 203.77 109.625 203.97 110.355 ;
      RECT 203.93 0.52 204.19 1.5 ;
      RECT 204.59 109.625 204.79 110.355 ;
      RECT 204.795 0.52 205.055 8.085 ;
      RECT 205.085 109.625 205.285 110.355 ;
      RECT 205.46 0.52 205.72 2.255 ;
      RECT 206.325 0.17 207.095 0.43 ;
      RECT 206.835 0.17 207.095 11.38 ;
      RECT 206.325 0.17 206.585 17.1 ;
      RECT 205.585 109.625 205.785 110.355 ;
      RECT 206.085 109.625 206.285 110.355 ;
      RECT 206.58 109.625 206.78 110.355 ;
      RECT 207.4 109.625 207.6 110.355 ;
      RECT 207.895 109.625 208.095 110.355 ;
      RECT 208.395 109.625 208.595 110.355 ;
      RECT 208.895 109.625 209.095 110.355 ;
      RECT 209.39 109.625 209.59 110.355 ;
      RECT 210.21 109.625 210.41 110.355 ;
      RECT 210.705 109.625 210.905 110.355 ;
      RECT 211.205 109.625 211.405 110.355 ;
      RECT 211.705 109.625 211.905 110.355 ;
      RECT 212.2 109.625 212.4 110.355 ;
      RECT 213.02 109.625 213.22 110.355 ;
      RECT 213.515 109.625 213.715 110.355 ;
      RECT 214.015 109.625 214.215 110.355 ;
      RECT 214.515 109.625 214.715 110.355 ;
      RECT 216.055 0.17 216.825 0.43 ;
      RECT 216.055 0.17 216.315 13.055 ;
      RECT 216.565 0.17 216.825 13.055 ;
      RECT 215.01 109.625 215.21 110.355 ;
      RECT 215.83 109.625 216.03 110.355 ;
      RECT 216.325 109.625 216.525 110.355 ;
      RECT 216.825 109.625 217.025 110.355 ;
      RECT 217.325 109.625 217.525 110.355 ;
      RECT 217.82 109.625 218.02 110.355 ;
      RECT 218.64 109.625 218.84 110.355 ;
      RECT 219.775 0.8 220.545 1.57 ;
      RECT 219.775 0.3 220.035 13.03 ;
      RECT 220.285 0.3 220.545 13.03 ;
      RECT 219.135 109.625 219.335 110.355 ;
      RECT 219.635 109.625 219.835 110.355 ;
      RECT 220.135 109.625 220.335 110.355 ;
      RECT 220.63 109.625 220.83 110.355 ;
      RECT 221 0.52 221.26 2.255 ;
      RECT 221.45 109.625 221.65 110.355 ;
      RECT 221.945 109.625 222.145 110.355 ;
      RECT 222.445 109.625 222.645 110.355 ;
      RECT 222.53 0.52 222.79 2.255 ;
      RECT 222.945 109.625 223.145 110.355 ;
      RECT 223.44 109.625 223.64 110.355 ;
      RECT 224.26 109.625 224.46 110.355 ;
      RECT 224.755 109.625 224.955 110.355 ;
      RECT 225.255 109.625 225.455 110.355 ;
      RECT 225.755 109.625 225.955 110.355 ;
      RECT 226.25 109.625 226.45 110.355 ;
      RECT 226.41 0.52 226.67 1.5 ;
      RECT 227.07 109.625 227.27 110.355 ;
      RECT 227.275 0.52 227.535 8.085 ;
      RECT 227.565 109.625 227.765 110.355 ;
      RECT 227.94 0.52 228.2 2.255 ;
      RECT 228.805 0.17 229.575 0.43 ;
      RECT 229.315 0.17 229.575 11.38 ;
      RECT 228.805 0.17 229.065 17.1 ;
      RECT 228.065 109.625 228.265 110.355 ;
      RECT 228.565 109.625 228.765 110.355 ;
      RECT 229.06 109.625 229.26 110.355 ;
      RECT 229.88 109.625 230.08 110.355 ;
      RECT 230.375 109.625 230.575 110.355 ;
      RECT 230.875 109.625 231.075 110.355 ;
      RECT 231.375 109.625 231.575 110.355 ;
      RECT 231.87 109.625 232.07 110.355 ;
      RECT 232.69 109.625 232.89 110.355 ;
      RECT 233.185 109.625 233.385 110.355 ;
      RECT 233.685 109.625 233.885 110.355 ;
      RECT 234.185 109.625 234.385 110.355 ;
      RECT 234.68 109.625 234.88 110.355 ;
      RECT 235.5 109.625 235.7 110.355 ;
      RECT 236.495 37.065 236.695 110.355 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 0 0.52 236.8 110.38 ;
      RECT 228.46 0 236.8 110.38 ;
      RECT 223.05 0 226.15 110.38 ;
      RECT 221.52 0 222.27 110.38 ;
      RECT 205.98 0 220.74 110.38 ;
      RECT 200.57 0 203.67 110.38 ;
      RECT 199.04 0 199.79 110.38 ;
      RECT 183.5 0 198.26 110.38 ;
      RECT 178.09 0 181.19 110.38 ;
      RECT 176.56 0 177.31 110.38 ;
      RECT 161.02 0 175.78 110.38 ;
      RECT 155.61 0 158.71 110.38 ;
      RECT 154.08 0 154.83 110.38 ;
      RECT 135 0.17 153.3 110.38 ;
      RECT 135.01 0 153.3 110.38 ;
      RECT 125.31 0 134.23 110.38 ;
      RECT 119.71 0 120.97 110.38 ;
      RECT 118.18 0 118.42 110.38 ;
      RECT 116.65 0 116.89 110.38 ;
      RECT 113.59 0 113.83 110.38 ;
      RECT 112.06 0 112.3 110.38 ;
      RECT 104.4 0 110.77 110.38 ;
      RECT 101.85 0 102.11 110.38 ;
      RECT 100.33 0 101.08 110.38 ;
      RECT 83.5 0 99.56 110.38 ;
      RECT 81.97 0 82.72 110.38 ;
      RECT 78.09 0 81.19 110.38 ;
      RECT 61.02 0 75.78 110.38 ;
      RECT 59.49 0 60.24 110.38 ;
      RECT 55.61 0 58.71 110.38 ;
      RECT 38.54 0 53.3 110.38 ;
      RECT 37.01 0 37.76 110.38 ;
      RECT 33.13 0 36.23 110.38 ;
      RECT 16.06 0 30.82 110.38 ;
      RECT 14.53 0 15.28 110.38 ;
      RECT 10.65 0 13.75 110.38 ;
      RECT 0 0 8.34 110.38 ;
    LAYER Metal3 ;
      RECT 0 0 236.8 110.38 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 138.09 0 145.17 110.38 ;
      RECT 132.94 0 134.76 110.38 ;
      RECT 127.79 0 129.61 110.38 ;
      RECT 232.8 0 236.8 110.38 ;
      RECT 227.18 0 229.47 110.38 ;
      RECT 227.18 30.685 236.8 36.805 ;
      RECT 221.56 0 223.85 110.38 ;
      RECT 215.94 0 218.23 110.38 ;
      RECT 215.94 30.685 223.85 36.805 ;
      RECT 210.32 0 212.61 110.38 ;
      RECT 204.7 0 206.99 110.38 ;
      RECT 204.7 30.685 212.61 36.805 ;
      RECT 199.08 0 201.37 110.38 ;
      RECT 193.46 0 195.75 110.38 ;
      RECT 193.46 30.685 201.37 36.805 ;
      RECT 187.84 0 190.13 110.38 ;
      RECT 46.67 30.685 54.58 36.805 ;
      RECT 41.05 0 43.34 110.38 ;
      RECT 35.43 0 37.72 110.38 ;
      RECT 35.43 30.685 43.34 36.805 ;
      RECT 29.81 0 32.1 110.38 ;
      RECT 24.19 0 26.48 110.38 ;
      RECT 24.19 30.685 32.1 36.805 ;
      RECT 18.57 0 20.86 110.38 ;
      RECT 12.95 0 15.24 110.38 ;
      RECT 12.95 30.685 20.86 36.805 ;
      RECT 7.33 0 9.62 110.38 ;
      RECT 0 0 4 110.38 ;
      RECT 0 30.685 9.62 36.805 ;
      RECT 182.22 0 184.51 110.38 ;
      RECT 182.22 30.685 190.13 36.805 ;
      RECT 176.6 0 178.89 110.38 ;
      RECT 170.98 0 173.27 110.38 ;
      RECT 170.98 30.685 178.89 36.805 ;
      RECT 165.36 0 167.65 110.38 ;
      RECT 159.74 0 162.03 110.38 ;
      RECT 159.74 30.685 167.65 36.805 ;
      RECT 154.12 0 156.41 110.38 ;
      RECT 148.5 0 150.79 110.38 ;
      RECT 148.5 30.685 156.41 36.805 ;
      RECT 122.64 0 124.46 110.38 ;
      RECT 117.49 0 119.31 110.38 ;
      RECT 112.34 0 114.16 110.38 ;
      RECT 107.19 0 109.01 110.38 ;
      RECT 102.04 0 103.86 110.38 ;
      RECT 91.63 0 98.71 110.38 ;
      RECT 86.01 0 88.3 110.38 ;
      RECT 80.39 0 82.68 110.38 ;
      RECT 80.39 30.685 88.3 36.805 ;
      RECT 74.77 0 77.06 110.38 ;
      RECT 69.15 0 71.44 110.38 ;
      RECT 69.15 30.685 77.06 36.805 ;
      RECT 63.53 0 65.82 110.38 ;
      RECT 57.91 0 60.2 110.38 ;
      RECT 57.91 30.685 65.82 36.805 ;
      RECT 52.29 0 54.58 110.38 ;
      RECT 46.67 0 48.96 110.38 ;
  END
END RM_IHPSG13_1P_512x8_c3_bm_bist

END LIBRARY
