# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Tue Sep  9 10:49:24 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_1024x16_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_1024x16_c2_bm_bist 0 0 ;
  SIZE 402.61 BY 385.37 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.71 0 266.97 0.26 ;
    END
  END A_DIN[8]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.64 0 135.9 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.22 0 267.48 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.13 0 135.39 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 275.38 0 275.64 0.26 ;
    END
  END A_BM[8]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.97 0 127.23 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 274.005 0 274.265 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 128.345 0 128.605 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.57 0 259.83 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.78 0 143.04 0.26 ;
    END
  END A_DOUT[7]
  PIN B_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 269.26 0 269.52 0.26 ;
    END
  END B_DIN[8]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.09 0 133.35 0.26 ;
    END
  END B_DIN[7]
  PIN B_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.73 0 267.99 0.26 ;
    END
  END B_BIST_DIN[8]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.62 0 134.88 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 260.745 0 261.005 0.26 ;
    END
  END B_BM[8]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 141.605 0 141.865 0.26 ;
    END
  END B_BM[7]
  PIN B_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 262.275 0 262.535 0.26 ;
    END
  END B_BIST_BM[8]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 140.075 0 140.335 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.4 0 276.66 0.26 ;
    END
  END B_DOUT[8]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.95 0 126.21 0.26 ;
    END
  END B_DOUT[7]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 383.205 0 387.625 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 365.525 0 369.945 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.845 0 352.265 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.165 0 334.585 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 312.485 0 316.905 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.805 0 299.225 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 277.125 0 281.545 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 259.445 0 263.865 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 238.525 0 241.335 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 228.225 0 231.035 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.775 0 215.585 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 202.475 0 205.285 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 197.325 0 200.135 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 187.025 0 189.835 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 171.575 0 174.385 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.275 0 164.085 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.745 0 143.165 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.065 0 125.485 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.385 0 107.805 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.705 0 90.125 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 385.37 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 392.045 0 396.465 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.365 0 378.785 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 356.685 0 361.105 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 339.005 0 343.425 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 321.325 0 325.745 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 303.645 0 308.065 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.965 0 290.385 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 268.285 0 272.705 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 233.375 0 236.185 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.075 0 225.885 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.925 0 220.735 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.625 0 210.435 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 192.175 0 194.985 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 181.875 0 184.685 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 176.725 0 179.535 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.425 0 169.235 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 0 134.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 0 116.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 0 98.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 0 81.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 392.045 53.41 396.465 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.365 53.41 378.785 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 356.685 53.41 361.105 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 339.005 53.41 343.425 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 321.325 53.41 325.745 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 303.645 53.41 308.065 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.965 53.41 290.385 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 268.285 53.41 272.705 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 53.41 134.325 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 53.41 116.645 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 53.41 98.965 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 53.41 81.285 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 385.37 ;
    END
  END VDDARRAY!
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.39 0 284.65 0.26 ;
    END
  END A_DIN[9]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.96 0 118.22 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.9 0 285.16 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.45 0 117.71 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.06 0 293.32 0.26 ;
    END
  END A_BM[9]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.29 0 109.55 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 291.685 0 291.945 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.665 0 110.925 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.25 0 277.51 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.1 0 125.36 0.26 ;
    END
  END A_DOUT[6]
  PIN B_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 286.94 0 287.2 0.26 ;
    END
  END B_DIN[9]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.41 0 115.67 0.26 ;
    END
  END B_DIN[6]
  PIN B_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 285.41 0 285.67 0.26 ;
    END
  END B_BIST_DIN[9]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.94 0 117.2 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 278.425 0 278.685 0.26 ;
    END
  END B_BM[9]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.925 0 124.185 0.26 ;
    END
  END B_BM[6]
  PIN B_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 279.955 0 280.215 0.26 ;
    END
  END B_BIST_BM[9]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.395 0 122.655 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.08 0 294.34 0.26 ;
    END
  END B_DOUT[9]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.27 0 108.53 0.26 ;
    END
  END B_DOUT[6]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 302.07 0 302.33 0.26 ;
    END
  END A_DIN[10]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.28 0 100.54 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 302.58 0 302.84 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.77 0 100.03 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 310.74 0 311 0.26 ;
    END
  END A_BM[10]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 91.61 0 91.87 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 309.365 0 309.625 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 92.985 0 93.245 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.93 0 295.19 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 107.42 0 107.68 0.26 ;
    END
  END A_DOUT[5]
  PIN B_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.62 0 304.88 0.26 ;
    END
  END B_DIN[10]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 97.73 0 97.99 0.26 ;
    END
  END B_DIN[5]
  PIN B_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 303.09 0 303.35 0.26 ;
    END
  END B_BIST_DIN[10]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.26 0 99.52 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 296.105 0 296.365 0.26 ;
    END
  END B_BM[10]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 106.245 0 106.505 0.26 ;
    END
  END B_BM[5]
  PIN B_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 297.635 0 297.895 0.26 ;
    END
  END B_BIST_BM[10]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.715 0 104.975 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.76 0 312.02 0.26 ;
    END
  END B_DOUT[10]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 90.59 0 90.85 0.26 ;
    END
  END B_DOUT[5]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 319.75 0 320.01 0.26 ;
    END
  END A_DIN[11]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.6 0 82.86 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 320.26 0 320.52 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.09 0 82.35 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 328.42 0 328.68 0.26 ;
    END
  END A_BM[11]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 73.93 0 74.19 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.045 0 327.305 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 75.305 0 75.565 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 312.61 0 312.87 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.74 0 90 0.26 ;
    END
  END A_DOUT[4]
  PIN B_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 322.3 0 322.56 0.26 ;
    END
  END B_DIN[11]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 80.05 0 80.31 0.26 ;
    END
  END B_DIN[4]
  PIN B_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 320.77 0 321.03 0.26 ;
    END
  END B_BIST_DIN[11]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.58 0 81.84 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 313.785 0 314.045 0.26 ;
    END
  END B_BM[11]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.565 0 88.825 0.26 ;
    END
  END B_BM[4]
  PIN B_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.315 0 315.575 0.26 ;
    END
  END B_BIST_BM[11]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 87.035 0 87.295 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 329.44 0 329.7 0.26 ;
    END
  END B_DOUT[11]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.91 0 73.17 0.26 ;
    END
  END B_DOUT[4]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.43 0 337.69 0.26 ;
    END
  END A_DIN[12]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.94 0 338.2 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.1 0 346.36 0.26 ;
    END
  END A_BM[12]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 344.725 0 344.985 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 330.29 0 330.55 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.98 0 340.24 0.26 ;
    END
  END B_DIN[12]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.45 0 338.71 0.26 ;
    END
  END B_BIST_DIN[12]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 331.465 0 331.725 0.26 ;
    END
  END B_BM[12]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 332.995 0 333.255 0.26 ;
    END
  END B_BIST_BM[12]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.12 0 347.38 0.26 ;
    END
  END B_DOUT[12]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.11 0 355.37 0.26 ;
    END
  END A_DIN[13]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.62 0 355.88 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 363.78 0 364.04 0.26 ;
    END
  END A_BM[13]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.405 0 362.665 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.97 0 348.23 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 357.66 0 357.92 0.26 ;
    END
  END B_DIN[13]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.13 0 356.39 0.26 ;
    END
  END B_BIST_DIN[13]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.145 0 349.405 0.26 ;
    END
  END B_BM[13]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 350.675 0 350.935 0.26 ;
    END
  END B_BIST_BM[13]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.8 0 365.06 0.26 ;
    END
  END B_DOUT[13]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.79 0 373.05 0.26 ;
    END
  END A_DIN[14]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.3 0 373.56 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 381.46 0 381.72 0.26 ;
    END
  END A_BM[14]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 380.085 0 380.345 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 365.65 0 365.91 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 375.34 0 375.6 0.26 ;
    END
  END B_DIN[14]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.81 0 374.07 0.26 ;
    END
  END B_BIST_DIN[14]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 366.825 0 367.085 0.26 ;
    END
  END B_BM[14]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.355 0 368.615 0.26 ;
    END
  END B_BIST_BM[14]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.48 0 382.74 0.26 ;
    END
  END B_DOUT[14]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.47 0 390.73 0.26 ;
    END
  END A_DIN[15]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.98 0 391.24 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 399.14 0 399.4 0.26 ;
    END
  END A_BM[15]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 397.765 0 398.025 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 383.33 0 383.59 0.26 ;
    END
  END A_DOUT[15]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 393.02 0 393.28 0.26 ;
    END
  END B_DIN[15]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 391.49 0 391.75 0.26 ;
    END
  END B_BIST_DIN[15]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.505 0 384.765 0.26 ;
    END
  END B_BM[15]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 386.035 0 386.295 0.26 ;
    END
  END B_BIST_BM[15]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.16 0 400.42 0.26 ;
    END
  END B_DOUT[15]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.395 0 217.655 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.005 0 223.265 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 184.955 0 185.215 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.345 0 179.605 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.905 0 218.165 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.515 0 223.775 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 184.445 0 184.705 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.835 0 179.095 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 226.575 0 226.835 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 227.085 0 227.345 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 175.775 0 176.035 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 175.265 0 175.525 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 225.555 0 225.815 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 226.065 0 226.325 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 176.795 0 177.055 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 176.285 0 176.545 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.175 0 206.435 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.685 0 206.945 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.175 0 196.435 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.665 0 195.925 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.155 0 205.415 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.665 0 205.925 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 197.195 0 197.455 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.685 0 196.945 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 229.125 0 229.385 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.615 0 228.875 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 173.225 0 173.485 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 173.735 0 173.995 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.105 0 228.365 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.595 0 227.855 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 174.245 0 174.505 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 174.755 0 175.015 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.675 0 231.935 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.185 0 232.445 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN B_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 170.675 0 170.935 0.26 ;
    END
  END B_ADDR[8]
  PIN B_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 170.165 0 170.425 0.26 ;
    END
  END B_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 229.635 0 229.895 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 230.145 0 230.405 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN B_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.715 0 172.975 0.26 ;
    END
  END B_ADDR[9]
  PIN B_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.205 0 172.465 0.26 ;
    END
  END B_BIST_ADDR[9]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.865 0 216.125 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 219.435 0 219.695 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 218.925 0 219.185 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 216.375 0 216.635 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 236.775 0 237.035 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 186.485 0 186.745 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.915 0 183.175 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 183.425 0 183.685 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 185.975 0 186.235 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 165.575 0 165.835 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 146.7701 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 16.445 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.096283 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 218.415 0 218.675 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.335 0 214.595 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 220.965 0 221.225 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 220.455 0 220.715 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.845 0 215.105 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 147.2093 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 16.445 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.12299 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 183.935 0 184.195 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.015 0 188.275 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.385 0 181.645 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.895 0 182.155 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 187.505 0 187.765 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 402.61 385.37 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 385.34 ;
      RECT 1.135 384.61 1.335 385.34 ;
      RECT 1.545 384.61 1.905 385.34 ;
      RECT 2.115 384.61 2.315 385.34 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 384.61 2.97 385.34 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 384.61 3.54 385.34 ;
      RECT 3.835 384.61 4.035 385.34 ;
      RECT 4.33 384.61 4.69 385.34 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 384.61 5.1 385.34 ;
      RECT 5.555 384.61 5.755 385.34 ;
      RECT 5.965 384.61 6.325 385.34 ;
      RECT 6.535 384.61 6.735 385.34 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 384.61 7.39 385.34 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 384.61 7.96 385.34 ;
      RECT 8.255 384.61 8.455 385.34 ;
      RECT 8.75 384.61 9.11 385.34 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 384.61 9.52 385.34 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 384.61 10.175 385.34 ;
      RECT 10.385 384.61 10.745 385.34 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 384.61 11.155 385.34 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 384.61 11.81 385.34 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 384.61 12.38 385.34 ;
      RECT 12.675 384.61 12.875 385.34 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 384.61 13.53 385.34 ;
      RECT 13.74 384.61 13.94 385.34 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 384.61 14.595 385.34 ;
      RECT 14.805 384.61 15.165 385.34 ;
      RECT 15.375 384.61 15.575 385.34 ;
      RECT 16.03 384.61 16.23 385.34 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 384.61 16.8 385.34 ;
      RECT 17.095 384.61 17.295 385.34 ;
      RECT 17.59 384.61 17.95 385.34 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 384.61 18.36 385.34 ;
      RECT 18.815 384.61 19.015 385.34 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 384.61 19.585 385.34 ;
      RECT 19.795 384.61 19.995 385.34 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 384.61 20.65 385.34 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 384.61 21.22 385.34 ;
      RECT 21.515 384.61 21.715 385.34 ;
      RECT 22.01 384.61 22.37 385.34 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 384.61 22.78 385.34 ;
      RECT 23.235 384.61 23.435 385.34 ;
      RECT 23.645 384.61 24.005 385.34 ;
      RECT 24.215 384.61 24.415 385.34 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 384.61 25.07 385.34 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 384.61 25.64 385.34 ;
      RECT 25.935 384.61 26.135 385.34 ;
      RECT 26.43 384.61 26.79 385.34 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 384.61 27.2 385.34 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 384.61 27.855 385.34 ;
      RECT 28.065 384.61 28.425 385.34 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 384.61 28.835 385.34 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 384.61 29.49 385.34 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 384.61 30.06 385.34 ;
      RECT 30.355 384.61 30.555 385.34 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 384.61 31.21 385.34 ;
      RECT 31.42 384.61 31.62 385.34 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 384.61 32.275 385.34 ;
      RECT 32.485 384.61 32.845 385.34 ;
      RECT 33.055 384.61 33.255 385.34 ;
      RECT 33.71 384.61 33.91 385.34 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 384.61 34.48 385.34 ;
      RECT 34.775 384.61 34.975 385.34 ;
      RECT 35.27 384.61 35.63 385.34 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 384.61 36.04 385.34 ;
      RECT 36.495 384.61 36.695 385.34 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 384.61 37.265 385.34 ;
      RECT 37.475 384.61 37.675 385.34 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 384.61 38.33 385.34 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 384.61 38.9 385.34 ;
      RECT 39.195 384.61 39.395 385.34 ;
      RECT 39.69 384.61 40.05 385.34 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 384.61 40.46 385.34 ;
      RECT 40.915 384.61 41.115 385.34 ;
      RECT 41.325 384.61 41.685 385.34 ;
      RECT 41.895 384.61 42.095 385.34 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 384.61 42.75 385.34 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 384.61 43.32 385.34 ;
      RECT 43.615 384.61 43.815 385.34 ;
      RECT 44.11 384.61 44.47 385.34 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 384.61 44.88 385.34 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 384.61 45.535 385.34 ;
      RECT 45.745 384.61 46.105 385.34 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 384.61 46.515 385.34 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 384.61 47.17 385.34 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 384.61 47.74 385.34 ;
      RECT 48.035 384.61 48.235 385.34 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 384.61 48.89 385.34 ;
      RECT 49.1 384.61 49.3 385.34 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 384.61 49.955 385.34 ;
      RECT 50.165 384.61 50.525 385.34 ;
      RECT 50.735 384.61 50.935 385.34 ;
      RECT 51.39 384.61 51.59 385.34 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 384.61 52.16 385.34 ;
      RECT 52.455 384.61 52.655 385.34 ;
      RECT 52.95 384.61 53.31 385.34 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 384.61 53.72 385.34 ;
      RECT 54.175 384.61 54.375 385.34 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 384.61 54.945 385.34 ;
      RECT 55.155 384.61 55.355 385.34 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 384.61 56.01 385.34 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 384.61 56.58 385.34 ;
      RECT 56.875 384.61 57.075 385.34 ;
      RECT 57.37 384.61 57.73 385.34 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 384.61 58.14 385.34 ;
      RECT 58.595 384.61 58.795 385.34 ;
      RECT 59.005 384.61 59.365 385.34 ;
      RECT 59.575 384.61 59.775 385.34 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 384.61 60.43 385.34 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 384.61 61 385.34 ;
      RECT 61.295 384.61 61.495 385.34 ;
      RECT 61.79 384.61 62.15 385.34 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 384.61 62.56 385.34 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 384.61 63.215 385.34 ;
      RECT 63.425 384.61 63.785 385.34 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 384.61 64.195 385.34 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 384.61 64.85 385.34 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 384.61 65.42 385.34 ;
      RECT 65.715 384.61 65.915 385.34 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 384.61 66.57 385.34 ;
      RECT 66.78 384.61 66.98 385.34 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 384.61 67.635 385.34 ;
      RECT 67.845 384.61 68.205 385.34 ;
      RECT 68.415 384.61 68.615 385.34 ;
      RECT 69.07 384.61 69.27 385.34 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 384.61 69.84 385.34 ;
      RECT 70.135 384.61 70.335 385.34 ;
      RECT 70.63 384.61 70.99 385.34 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 384.61 71.4 385.34 ;
      RECT 71.855 384.61 72.055 385.34 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 72.265 384.61 72.625 385.34 ;
      RECT 72.835 384.61 73.035 385.34 ;
      RECT 72.91 0.52 73.17 7.78 ;
      RECT 73.42 0.3 73.68 5.235 ;
      RECT 73.49 384.61 73.69 385.34 ;
      RECT 73.93 0.52 74.19 5.57 ;
      RECT 73.9 384.61 74.26 385.34 ;
      RECT 74.555 384.61 74.755 385.34 ;
      RECT 75.05 384.61 75.41 385.34 ;
      RECT 75.305 0.52 75.565 6.28 ;
      RECT 75.62 384.61 75.82 385.34 ;
      RECT 76.275 384.61 76.475 385.34 ;
      RECT 76.685 384.61 77.045 385.34 ;
      RECT 77.255 384.61 77.455 385.34 ;
      RECT 76.99 0.18 77.76 0.88 ;
      RECT 77.91 384.61 78.11 385.34 ;
      RECT 78.01 0.3 78.27 8.7 ;
      RECT 78.32 384.61 78.68 385.34 ;
      RECT 78.975 384.61 79.175 385.34 ;
      RECT 79.47 384.61 79.83 385.34 ;
      RECT 80.56 0.155 81.33 0.445 ;
      RECT 80.56 0.155 80.82 8.665 ;
      RECT 81.07 0.155 81.33 8.665 ;
      RECT 80.04 384.61 80.24 385.34 ;
      RECT 80.05 0.52 80.31 9.955 ;
      RECT 80.695 384.61 80.895 385.34 ;
      RECT 81.105 384.61 81.465 385.34 ;
      RECT 81.58 0.52 81.84 11.315 ;
      RECT 81.675 384.61 81.875 385.34 ;
      RECT 82.09 0.52 82.35 13.45 ;
      RECT 82.33 384.61 82.53 385.34 ;
      RECT 82.6 0.52 82.86 14.115 ;
      RECT 82.74 384.61 83.1 385.34 ;
      RECT 83.395 384.61 83.595 385.34 ;
      RECT 84.795 0.155 85.565 0.445 ;
      RECT 84.795 0.155 85.055 13.21 ;
      RECT 85.305 0.155 85.565 13.21 ;
      RECT 83.89 384.61 84.25 385.34 ;
      RECT 84.46 384.61 84.66 385.34 ;
      RECT 85.815 0.18 86.585 0.88 ;
      RECT 85.815 0.18 86.075 12.9 ;
      RECT 86.325 0.18 86.585 12.9 ;
      RECT 85.115 384.61 85.315 385.34 ;
      RECT 85.525 384.61 85.885 385.34 ;
      RECT 86.095 384.61 86.295 385.34 ;
      RECT 86.75 384.61 86.95 385.34 ;
      RECT 87.035 0.52 87.295 2.82 ;
      RECT 87.16 384.61 87.52 385.34 ;
      RECT 87.815 384.61 88.015 385.34 ;
      RECT 88.31 384.61 88.67 385.34 ;
      RECT 88.565 0.52 88.825 2.82 ;
      RECT 88.88 384.61 89.08 385.34 ;
      RECT 89.535 384.61 89.735 385.34 ;
      RECT 89.74 0.52 90 4.315 ;
      RECT 89.945 384.61 90.305 385.34 ;
      RECT 90.515 384.61 90.715 385.34 ;
      RECT 90.59 0.52 90.85 7.78 ;
      RECT 91.1 0.3 91.36 5.235 ;
      RECT 91.17 384.61 91.37 385.34 ;
      RECT 91.61 0.52 91.87 5.57 ;
      RECT 91.58 384.61 91.94 385.34 ;
      RECT 92.235 384.61 92.435 385.34 ;
      RECT 92.73 384.61 93.09 385.34 ;
      RECT 92.985 0.52 93.245 6.28 ;
      RECT 93.3 384.61 93.5 385.34 ;
      RECT 93.955 384.61 94.155 385.34 ;
      RECT 94.365 384.61 94.725 385.34 ;
      RECT 94.935 384.61 95.135 385.34 ;
      RECT 94.67 0.18 95.44 0.88 ;
      RECT 95.59 384.61 95.79 385.34 ;
      RECT 95.69 0.3 95.95 8.7 ;
      RECT 96 384.61 96.36 385.34 ;
      RECT 96.655 384.61 96.855 385.34 ;
      RECT 97.15 384.61 97.51 385.34 ;
      RECT 98.24 0.155 99.01 0.445 ;
      RECT 98.24 0.155 98.5 8.665 ;
      RECT 98.75 0.155 99.01 8.665 ;
      RECT 97.72 384.61 97.92 385.34 ;
      RECT 97.73 0.52 97.99 9.955 ;
      RECT 98.375 384.61 98.575 385.34 ;
      RECT 98.785 384.61 99.145 385.34 ;
      RECT 99.26 0.52 99.52 11.315 ;
      RECT 99.355 384.61 99.555 385.34 ;
      RECT 99.77 0.52 100.03 13.45 ;
      RECT 100.01 384.61 100.21 385.34 ;
      RECT 100.28 0.52 100.54 14.115 ;
      RECT 100.42 384.61 100.78 385.34 ;
      RECT 101.075 384.61 101.275 385.34 ;
      RECT 102.475 0.155 103.245 0.445 ;
      RECT 102.475 0.155 102.735 13.21 ;
      RECT 102.985 0.155 103.245 13.21 ;
      RECT 101.57 384.61 101.93 385.34 ;
      RECT 102.14 384.61 102.34 385.34 ;
      RECT 103.495 0.18 104.265 0.88 ;
      RECT 103.495 0.18 103.755 12.9 ;
      RECT 104.005 0.18 104.265 12.9 ;
      RECT 102.795 384.61 102.995 385.34 ;
      RECT 103.205 384.61 103.565 385.34 ;
      RECT 103.775 384.61 103.975 385.34 ;
      RECT 104.43 384.61 104.63 385.34 ;
      RECT 104.715 0.52 104.975 2.82 ;
      RECT 104.84 384.61 105.2 385.34 ;
      RECT 105.495 384.61 105.695 385.34 ;
      RECT 105.99 384.61 106.35 385.34 ;
      RECT 106.245 0.52 106.505 2.82 ;
      RECT 106.56 384.61 106.76 385.34 ;
      RECT 107.215 384.61 107.415 385.34 ;
      RECT 107.42 0.52 107.68 4.315 ;
      RECT 107.625 384.61 107.985 385.34 ;
      RECT 108.195 384.61 108.395 385.34 ;
      RECT 108.27 0.52 108.53 7.78 ;
      RECT 108.78 0.3 109.04 5.235 ;
      RECT 108.85 384.61 109.05 385.34 ;
      RECT 109.29 0.52 109.55 5.57 ;
      RECT 109.26 384.61 109.62 385.34 ;
      RECT 109.915 384.61 110.115 385.34 ;
      RECT 110.41 384.61 110.77 385.34 ;
      RECT 110.665 0.52 110.925 6.28 ;
      RECT 110.98 384.61 111.18 385.34 ;
      RECT 111.635 384.61 111.835 385.34 ;
      RECT 112.045 384.61 112.405 385.34 ;
      RECT 112.615 384.61 112.815 385.34 ;
      RECT 112.35 0.18 113.12 0.88 ;
      RECT 113.27 384.61 113.47 385.34 ;
      RECT 113.37 0.3 113.63 8.7 ;
      RECT 113.68 384.61 114.04 385.34 ;
      RECT 114.335 384.61 114.535 385.34 ;
      RECT 114.83 384.61 115.19 385.34 ;
      RECT 115.92 0.155 116.69 0.445 ;
      RECT 115.92 0.155 116.18 8.665 ;
      RECT 116.43 0.155 116.69 8.665 ;
      RECT 115.4 384.61 115.6 385.34 ;
      RECT 115.41 0.52 115.67 9.955 ;
      RECT 116.055 384.61 116.255 385.34 ;
      RECT 116.465 384.61 116.825 385.34 ;
      RECT 116.94 0.52 117.2 11.315 ;
      RECT 117.035 384.61 117.235 385.34 ;
      RECT 117.45 0.52 117.71 13.45 ;
      RECT 117.69 384.61 117.89 385.34 ;
      RECT 117.96 0.52 118.22 14.115 ;
      RECT 118.1 384.61 118.46 385.34 ;
      RECT 118.755 384.61 118.955 385.34 ;
      RECT 120.155 0.155 120.925 0.445 ;
      RECT 120.155 0.155 120.415 13.21 ;
      RECT 120.665 0.155 120.925 13.21 ;
      RECT 119.25 384.61 119.61 385.34 ;
      RECT 119.82 384.61 120.02 385.34 ;
      RECT 121.175 0.18 121.945 0.88 ;
      RECT 121.175 0.18 121.435 12.9 ;
      RECT 121.685 0.18 121.945 12.9 ;
      RECT 120.475 384.61 120.675 385.34 ;
      RECT 120.885 384.61 121.245 385.34 ;
      RECT 121.455 384.61 121.655 385.34 ;
      RECT 122.11 384.61 122.31 385.34 ;
      RECT 122.395 0.52 122.655 2.82 ;
      RECT 122.52 384.61 122.88 385.34 ;
      RECT 123.175 384.61 123.375 385.34 ;
      RECT 123.67 384.61 124.03 385.34 ;
      RECT 123.925 0.52 124.185 2.82 ;
      RECT 124.24 384.61 124.44 385.34 ;
      RECT 124.895 384.61 125.095 385.34 ;
      RECT 125.1 0.52 125.36 4.315 ;
      RECT 125.305 384.61 125.665 385.34 ;
      RECT 125.875 384.61 126.075 385.34 ;
      RECT 125.95 0.52 126.21 7.78 ;
      RECT 126.46 0.3 126.72 5.235 ;
      RECT 126.53 384.61 126.73 385.34 ;
      RECT 126.97 0.52 127.23 5.57 ;
      RECT 126.94 384.61 127.3 385.34 ;
      RECT 127.595 384.61 127.795 385.34 ;
      RECT 128.09 384.61 128.45 385.34 ;
      RECT 128.345 0.52 128.605 6.28 ;
      RECT 128.66 384.61 128.86 385.34 ;
      RECT 129.315 384.61 129.515 385.34 ;
      RECT 129.725 384.61 130.085 385.34 ;
      RECT 130.295 384.61 130.495 385.34 ;
      RECT 130.03 0.18 130.8 0.88 ;
      RECT 130.95 384.61 131.15 385.34 ;
      RECT 131.05 0.3 131.31 8.7 ;
      RECT 131.36 384.61 131.72 385.34 ;
      RECT 132.015 384.61 132.215 385.34 ;
      RECT 132.51 384.61 132.87 385.34 ;
      RECT 133.6 0.155 134.37 0.445 ;
      RECT 133.6 0.155 133.86 8.665 ;
      RECT 134.11 0.155 134.37 8.665 ;
      RECT 133.08 384.61 133.28 385.34 ;
      RECT 133.09 0.52 133.35 9.955 ;
      RECT 133.735 384.61 133.935 385.34 ;
      RECT 134.145 384.61 134.505 385.34 ;
      RECT 134.62 0.52 134.88 11.315 ;
      RECT 134.715 384.61 134.915 385.34 ;
      RECT 135.13 0.52 135.39 13.45 ;
      RECT 135.37 384.61 135.57 385.34 ;
      RECT 135.64 0.52 135.9 14.115 ;
      RECT 135.78 384.61 136.14 385.34 ;
      RECT 136.435 384.61 136.635 385.34 ;
      RECT 137.835 0.155 138.605 0.445 ;
      RECT 137.835 0.155 138.095 13.21 ;
      RECT 138.345 0.155 138.605 13.21 ;
      RECT 136.93 384.61 137.29 385.34 ;
      RECT 137.5 384.61 137.7 385.34 ;
      RECT 138.855 0.18 139.625 0.88 ;
      RECT 138.855 0.18 139.115 12.9 ;
      RECT 139.365 0.18 139.625 12.9 ;
      RECT 138.155 384.61 138.355 385.34 ;
      RECT 138.565 384.61 138.925 385.34 ;
      RECT 139.135 384.61 139.335 385.34 ;
      RECT 139.79 384.61 139.99 385.34 ;
      RECT 140.075 0.52 140.335 2.82 ;
      RECT 140.2 384.61 140.56 385.34 ;
      RECT 140.855 384.61 141.055 385.34 ;
      RECT 141.35 384.61 141.71 385.34 ;
      RECT 141.605 0.52 141.865 2.82 ;
      RECT 141.92 384.61 142.12 385.34 ;
      RECT 142.575 384.61 142.775 385.34 ;
      RECT 143.8 0.17 144.57 0.43 ;
      RECT 143.8 0.17 144.06 8.7 ;
      RECT 144.31 0.17 144.57 8.7 ;
      RECT 142.78 0.52 143.04 4.315 ;
      RECT 144.82 0.18 145.59 0.88 ;
      RECT 144.82 0.18 145.08 8.7 ;
      RECT 145.33 0.18 145.59 8.7 ;
      RECT 145.84 0.17 146.61 0.43 ;
      RECT 145.84 0.17 146.1 8.7 ;
      RECT 146.35 0.17 146.61 8.7 ;
      RECT 146.86 0.18 147.63 0.88 ;
      RECT 146.86 0.18 147.12 8.7 ;
      RECT 147.37 0.18 147.63 8.7 ;
      RECT 147.88 0.17 148.65 0.43 ;
      RECT 147.88 0.17 148.14 8.7 ;
      RECT 148.39 0.17 148.65 8.7 ;
      RECT 148.9 0.18 149.67 0.88 ;
      RECT 148.9 0.18 149.16 8.7 ;
      RECT 149.41 0.18 149.67 8.7 ;
      RECT 149.92 0.17 150.69 0.43 ;
      RECT 149.92 0.17 150.18 8.7 ;
      RECT 150.43 0.17 150.69 8.7 ;
      RECT 150.94 0.18 151.71 0.88 ;
      RECT 150.94 0.18 151.2 8.7 ;
      RECT 151.45 0.18 151.71 8.7 ;
      RECT 151.96 0.17 152.73 0.43 ;
      RECT 151.96 0.17 152.22 8.7 ;
      RECT 152.47 0.17 152.73 8.7 ;
      RECT 152.98 0.18 153.75 0.88 ;
      RECT 152.98 0.18 153.24 8.7 ;
      RECT 153.49 0.18 153.75 8.7 ;
      RECT 154 0.17 154.77 0.43 ;
      RECT 154 0.17 154.26 8.7 ;
      RECT 154.51 0.17 154.77 8.7 ;
      RECT 155.02 0.18 155.79 0.88 ;
      RECT 155.02 0.18 155.28 8.7 ;
      RECT 155.53 0.18 155.79 8.7 ;
      RECT 156.04 0.17 156.81 0.43 ;
      RECT 156.04 0.17 156.3 8.7 ;
      RECT 156.55 0.17 156.81 8.7 ;
      RECT 157.06 0.18 157.83 0.88 ;
      RECT 157.06 0.18 157.32 8.7 ;
      RECT 157.57 0.18 157.83 8.7 ;
      RECT 158.08 0.17 158.85 0.43 ;
      RECT 158.08 0.17 158.34 8.7 ;
      RECT 158.59 0.17 158.85 8.7 ;
      RECT 159.1 0.18 159.87 0.88 ;
      RECT 159.1 0.18 159.36 8.7 ;
      RECT 159.61 0.18 159.87 8.7 ;
      RECT 142.985 384.61 143.345 385.34 ;
      RECT 143.555 384.61 143.755 385.34 ;
      RECT 161.495 0.18 162.265 0.88 ;
      RECT 161.495 0.18 161.755 8.7 ;
      RECT 162.005 0.18 162.265 8.7 ;
      RECT 162.515 0.17 163.285 0.43 ;
      RECT 162.515 0.17 162.775 8.7 ;
      RECT 163.025 0.17 163.285 8.7 ;
      RECT 144.38 384.53 144.58 385.34 ;
      RECT 160.475 0.3 160.735 8.7 ;
      RECT 164.555 0.18 165.325 0.88 ;
      RECT 164.555 0.18 164.815 8.7 ;
      RECT 165.065 0.18 165.325 8.7 ;
      RECT 160.985 0.3 161.245 8.7 ;
      RECT 163.535 0 163.795 8.7 ;
      RECT 164.045 0 164.305 8.7 ;
      RECT 165.575 0.52 165.835 8.7 ;
      RECT 166.085 0.3 166.345 8.7 ;
      RECT 166.595 0.3 166.855 8.7 ;
      RECT 167.105 0.3 167.365 8.7 ;
      RECT 167.615 0.3 167.875 8.7 ;
      RECT 168.125 0.3 168.385 8.7 ;
      RECT 168.635 0.3 168.895 8.7 ;
      RECT 169.145 0.3 169.405 8.7 ;
      RECT 171.185 0.18 171.955 0.88 ;
      RECT 171.185 0.18 171.445 8.7 ;
      RECT 171.695 0.18 171.955 8.7 ;
      RECT 169.655 0.3 169.915 8.7 ;
      RECT 170.165 0.52 170.425 8.7 ;
      RECT 170.675 0.52 170.935 8.7 ;
      RECT 172.205 0.52 172.465 8.7 ;
      RECT 172.715 0.52 172.975 8.7 ;
      RECT 173.225 0.52 173.485 8.7 ;
      RECT 173.735 0.52 173.995 8.7 ;
      RECT 174.245 0.52 174.505 8.7 ;
      RECT 174.755 0.52 175.015 8.7 ;
      RECT 175.265 0.52 175.525 8.7 ;
      RECT 175.775 0.52 176.035 8.7 ;
      RECT 176.285 0.52 176.545 8.7 ;
      RECT 176.795 0.52 177.055 8.7 ;
      RECT 177.305 0.3 177.565 8.7 ;
      RECT 177.815 0.3 178.075 8.7 ;
      RECT 178.325 0.3 178.585 8.7 ;
      RECT 178.835 0.52 179.095 8.7 ;
      RECT 179.345 0.52 179.605 8.7 ;
      RECT 179.855 0.3 180.115 8.7 ;
      RECT 180.365 0.3 180.625 8.7 ;
      RECT 180.875 0.3 181.135 8.7 ;
      RECT 181.385 0.52 181.645 8.7 ;
      RECT 181.895 0.52 182.155 8.7 ;
      RECT 182.405 0.3 182.665 8.7 ;
      RECT 182.915 0.52 183.175 8.7 ;
      RECT 183.425 0.52 183.685 8.7 ;
      RECT 183.935 0.52 184.195 8.7 ;
      RECT 184.445 0.52 184.705 8.7 ;
      RECT 184.955 0.52 185.215 8.7 ;
      RECT 185.465 0.3 185.725 8.7 ;
      RECT 185.975 0.52 186.235 8.7 ;
      RECT 186.485 0.52 186.745 8.7 ;
      RECT 186.995 0.3 187.255 8.7 ;
      RECT 187.505 0.52 187.765 8.7 ;
      RECT 189.545 0.17 190.315 0.43 ;
      RECT 189.545 0.17 189.805 8.7 ;
      RECT 190.055 0.17 190.315 8.7 ;
      RECT 188.015 0.52 188.275 8.7 ;
      RECT 188.525 0.3 188.785 8.7 ;
      RECT 189.035 0.3 189.295 8.7 ;
      RECT 192.095 0.17 192.865 0.43 ;
      RECT 192.095 0.17 192.355 8.7 ;
      RECT 192.605 0.17 192.865 8.7 ;
      RECT 190.565 0.3 190.825 8.7 ;
      RECT 193.625 0.18 194.395 0.88 ;
      RECT 193.625 0.18 193.885 8.7 ;
      RECT 194.135 0.18 194.395 8.7 ;
      RECT 191.075 0.3 191.335 8.7 ;
      RECT 191.585 0.3 191.845 8.7 ;
      RECT 193.115 0.3 193.375 8.7 ;
      RECT 194.645 0 194.905 8.7 ;
      RECT 195.155 0 195.415 8.7 ;
      RECT 195.665 0.52 195.925 8.7 ;
      RECT 196.175 0.52 196.435 8.7 ;
      RECT 196.685 0.52 196.945 8.7 ;
      RECT 197.195 0.52 197.455 8.7 ;
      RECT 197.705 0 197.965 8.7 ;
      RECT 198.215 0 198.475 8.7 ;
      RECT 198.725 0.3 198.985 8.7 ;
      RECT 199.235 0.3 199.495 8.7 ;
      RECT 199.745 0 200.005 8.7 ;
      RECT 200.255 0 200.515 8.7 ;
      RECT 200.765 0.3 201.025 8.7 ;
      RECT 201.585 0.3 201.845 8.7 ;
      RECT 202.095 0 202.355 8.7 ;
      RECT 202.605 0 202.865 8.7 ;
      RECT 203.115 0.3 203.375 8.7 ;
      RECT 203.625 0.3 203.885 8.7 ;
      RECT 204.135 0 204.395 8.7 ;
      RECT 204.645 0 204.905 8.7 ;
      RECT 205.155 0.52 205.415 8.7 ;
      RECT 205.665 0.52 205.925 8.7 ;
      RECT 206.175 0.52 206.435 8.7 ;
      RECT 208.215 0.18 208.985 0.88 ;
      RECT 208.215 0.18 208.475 8.7 ;
      RECT 208.725 0.18 208.985 8.7 ;
      RECT 206.685 0.52 206.945 8.7 ;
      RECT 209.745 0.17 210.515 0.43 ;
      RECT 209.745 0.17 210.005 8.7 ;
      RECT 210.255 0.17 210.515 8.7 ;
      RECT 207.195 0 207.455 8.7 ;
      RECT 207.705 0 207.965 8.7 ;
      RECT 209.235 0.3 209.495 8.7 ;
      RECT 212.295 0.17 213.065 0.43 ;
      RECT 212.295 0.17 212.555 8.7 ;
      RECT 212.805 0.17 213.065 8.7 ;
      RECT 210.765 0.3 211.025 8.7 ;
      RECT 211.275 0.3 211.535 8.7 ;
      RECT 211.785 0.3 212.045 8.7 ;
      RECT 213.315 0.3 213.575 8.7 ;
      RECT 213.825 0.3 214.085 8.7 ;
      RECT 214.335 0.52 214.595 8.7 ;
      RECT 214.845 0.52 215.105 8.7 ;
      RECT 215.355 0.3 215.615 8.7 ;
      RECT 215.865 0.52 216.125 8.7 ;
      RECT 216.375 0.52 216.635 8.7 ;
      RECT 216.885 0.3 217.145 8.7 ;
      RECT 217.395 0.52 217.655 8.7 ;
      RECT 217.905 0.52 218.165 8.7 ;
      RECT 218.415 0.52 218.675 8.7 ;
      RECT 218.925 0.52 219.185 8.7 ;
      RECT 219.435 0.52 219.695 8.7 ;
      RECT 219.945 0.3 220.205 8.7 ;
      RECT 220.455 0.52 220.715 8.7 ;
      RECT 220.965 0.52 221.225 8.7 ;
      RECT 221.475 0.3 221.735 8.7 ;
      RECT 221.985 0.3 222.245 8.7 ;
      RECT 222.495 0.3 222.755 8.7 ;
      RECT 223.005 0.52 223.265 8.7 ;
      RECT 223.515 0.52 223.775 8.7 ;
      RECT 224.025 0.3 224.285 8.7 ;
      RECT 224.535 0.3 224.795 8.7 ;
      RECT 225.045 0.3 225.305 8.7 ;
      RECT 225.555 0.52 225.815 8.7 ;
      RECT 226.065 0.52 226.325 8.7 ;
      RECT 226.575 0.52 226.835 8.7 ;
      RECT 227.085 0.52 227.345 8.7 ;
      RECT 227.595 0.52 227.855 8.7 ;
      RECT 228.105 0.52 228.365 8.7 ;
      RECT 228.615 0.52 228.875 8.7 ;
      RECT 230.655 0.18 231.425 0.88 ;
      RECT 230.655 0.18 230.915 8.7 ;
      RECT 231.165 0.18 231.425 8.7 ;
      RECT 229.125 0.52 229.385 8.7 ;
      RECT 229.635 0.52 229.895 8.7 ;
      RECT 230.145 0.52 230.405 8.7 ;
      RECT 231.675 0.52 231.935 8.7 ;
      RECT 232.185 0.52 232.445 8.7 ;
      RECT 232.695 0.3 232.955 8.7 ;
      RECT 233.205 0.3 233.465 8.7 ;
      RECT 233.715 0.3 233.975 8.7 ;
      RECT 234.225 0.3 234.485 8.7 ;
      RECT 234.735 0.3 234.995 8.7 ;
      RECT 235.245 0.3 235.505 8.7 ;
      RECT 237.285 0.18 238.055 0.88 ;
      RECT 237.285 0.18 237.545 8.7 ;
      RECT 237.795 0.18 238.055 8.7 ;
      RECT 235.755 0.3 236.015 8.7 ;
      RECT 236.265 0.3 236.525 8.7 ;
      RECT 239.325 0.17 240.095 0.43 ;
      RECT 239.325 0.17 239.585 8.7 ;
      RECT 239.835 0.17 240.095 8.7 ;
      RECT 240.345 0.18 241.115 0.88 ;
      RECT 240.345 0.18 240.605 8.7 ;
      RECT 240.855 0.18 241.115 8.7 ;
      RECT 236.775 0.52 237.035 8.7 ;
      RECT 238.305 0 238.565 8.7 ;
      RECT 242.74 0.18 243.51 0.88 ;
      RECT 242.74 0.18 243 8.7 ;
      RECT 243.25 0.18 243.51 8.7 ;
      RECT 243.76 0.17 244.53 0.43 ;
      RECT 243.76 0.17 244.02 8.7 ;
      RECT 244.27 0.17 244.53 8.7 ;
      RECT 244.78 0.18 245.55 0.88 ;
      RECT 244.78 0.18 245.04 8.7 ;
      RECT 245.29 0.18 245.55 8.7 ;
      RECT 245.8 0.17 246.57 0.43 ;
      RECT 245.8 0.17 246.06 8.7 ;
      RECT 246.31 0.17 246.57 8.7 ;
      RECT 246.82 0.18 247.59 0.88 ;
      RECT 246.82 0.18 247.08 8.7 ;
      RECT 247.33 0.18 247.59 8.7 ;
      RECT 247.84 0.17 248.61 0.43 ;
      RECT 247.84 0.17 248.1 8.7 ;
      RECT 248.35 0.17 248.61 8.7 ;
      RECT 248.86 0.18 249.63 0.88 ;
      RECT 248.86 0.18 249.12 8.7 ;
      RECT 249.37 0.18 249.63 8.7 ;
      RECT 249.88 0.17 250.65 0.43 ;
      RECT 249.88 0.17 250.14 8.7 ;
      RECT 250.39 0.17 250.65 8.7 ;
      RECT 250.9 0.18 251.67 0.88 ;
      RECT 250.9 0.18 251.16 8.7 ;
      RECT 251.41 0.18 251.67 8.7 ;
      RECT 251.92 0.17 252.69 0.43 ;
      RECT 251.92 0.17 252.18 8.7 ;
      RECT 252.43 0.17 252.69 8.7 ;
      RECT 252.94 0.18 253.71 0.88 ;
      RECT 252.94 0.18 253.2 8.7 ;
      RECT 253.45 0.18 253.71 8.7 ;
      RECT 253.96 0.17 254.73 0.43 ;
      RECT 253.96 0.17 254.22 8.7 ;
      RECT 254.47 0.17 254.73 8.7 ;
      RECT 254.98 0.18 255.75 0.88 ;
      RECT 254.98 0.18 255.24 8.7 ;
      RECT 255.49 0.18 255.75 8.7 ;
      RECT 256 0.17 256.77 0.43 ;
      RECT 256 0.17 256.26 8.7 ;
      RECT 256.51 0.17 256.77 8.7 ;
      RECT 257.02 0.18 257.79 0.88 ;
      RECT 257.02 0.18 257.28 8.7 ;
      RECT 257.53 0.18 257.79 8.7 ;
      RECT 238.815 0 239.075 8.7 ;
      RECT 258.04 0.17 258.81 0.43 ;
      RECT 258.04 0.17 258.3 8.7 ;
      RECT 258.55 0.17 258.81 8.7 ;
      RECT 241.365 0.3 241.625 8.7 ;
      RECT 241.875 0.3 242.135 8.7 ;
      RECT 258.03 384.53 258.23 385.34 ;
      RECT 258.855 384.61 259.055 385.34 ;
      RECT 259.265 384.61 259.625 385.34 ;
      RECT 259.57 0.52 259.83 4.315 ;
      RECT 259.835 384.61 260.035 385.34 ;
      RECT 260.49 384.61 260.69 385.34 ;
      RECT 260.745 0.52 261.005 2.82 ;
      RECT 260.9 384.61 261.26 385.34 ;
      RECT 261.555 384.61 261.755 385.34 ;
      RECT 262.05 384.61 262.41 385.34 ;
      RECT 262.985 0.18 263.755 0.88 ;
      RECT 262.985 0.18 263.245 12.9 ;
      RECT 263.495 0.18 263.755 12.9 ;
      RECT 262.275 0.52 262.535 2.82 ;
      RECT 262.62 384.61 262.82 385.34 ;
      RECT 264.005 0.155 264.775 0.445 ;
      RECT 264.005 0.155 264.265 13.21 ;
      RECT 264.515 0.155 264.775 13.21 ;
      RECT 263.275 384.61 263.475 385.34 ;
      RECT 263.685 384.61 264.045 385.34 ;
      RECT 264.255 384.61 264.455 385.34 ;
      RECT 264.91 384.61 265.11 385.34 ;
      RECT 265.32 384.61 265.68 385.34 ;
      RECT 265.975 384.61 266.175 385.34 ;
      RECT 266.47 384.61 266.83 385.34 ;
      RECT 266.71 0.52 266.97 14.115 ;
      RECT 267.04 384.61 267.24 385.34 ;
      RECT 267.22 0.52 267.48 13.45 ;
      RECT 267.695 384.61 267.895 385.34 ;
      RECT 268.24 0.155 269.01 0.445 ;
      RECT 268.24 0.155 268.5 8.665 ;
      RECT 268.75 0.155 269.01 8.665 ;
      RECT 267.73 0.52 267.99 11.315 ;
      RECT 268.105 384.61 268.465 385.34 ;
      RECT 268.675 384.61 268.875 385.34 ;
      RECT 269.26 0.52 269.52 9.955 ;
      RECT 269.33 384.61 269.53 385.34 ;
      RECT 269.74 384.61 270.1 385.34 ;
      RECT 270.395 384.61 270.595 385.34 ;
      RECT 270.89 384.61 271.25 385.34 ;
      RECT 271.3 0.3 271.56 8.7 ;
      RECT 271.46 384.61 271.66 385.34 ;
      RECT 272.115 384.61 272.315 385.34 ;
      RECT 271.81 0.18 272.58 0.88 ;
      RECT 272.525 384.61 272.885 385.34 ;
      RECT 273.095 384.61 273.295 385.34 ;
      RECT 273.75 384.61 273.95 385.34 ;
      RECT 274.005 0.52 274.265 6.28 ;
      RECT 274.16 384.61 274.52 385.34 ;
      RECT 274.815 384.61 275.015 385.34 ;
      RECT 275.38 0.52 275.64 5.57 ;
      RECT 275.31 384.61 275.67 385.34 ;
      RECT 275.88 384.61 276.08 385.34 ;
      RECT 275.89 0.3 276.15 5.235 ;
      RECT 276.4 0.52 276.66 7.78 ;
      RECT 276.535 384.61 276.735 385.34 ;
      RECT 276.945 384.61 277.305 385.34 ;
      RECT 277.25 0.52 277.51 4.315 ;
      RECT 277.515 384.61 277.715 385.34 ;
      RECT 278.17 384.61 278.37 385.34 ;
      RECT 278.425 0.52 278.685 2.82 ;
      RECT 278.58 384.61 278.94 385.34 ;
      RECT 279.235 384.61 279.435 385.34 ;
      RECT 279.73 384.61 280.09 385.34 ;
      RECT 280.665 0.18 281.435 0.88 ;
      RECT 280.665 0.18 280.925 12.9 ;
      RECT 281.175 0.18 281.435 12.9 ;
      RECT 279.955 0.52 280.215 2.82 ;
      RECT 280.3 384.61 280.5 385.34 ;
      RECT 281.685 0.155 282.455 0.445 ;
      RECT 281.685 0.155 281.945 13.21 ;
      RECT 282.195 0.155 282.455 13.21 ;
      RECT 280.955 384.61 281.155 385.34 ;
      RECT 281.365 384.61 281.725 385.34 ;
      RECT 281.935 384.61 282.135 385.34 ;
      RECT 282.59 384.61 282.79 385.34 ;
      RECT 283 384.61 283.36 385.34 ;
      RECT 283.655 384.61 283.855 385.34 ;
      RECT 284.15 384.61 284.51 385.34 ;
      RECT 284.39 0.52 284.65 14.115 ;
      RECT 284.72 384.61 284.92 385.34 ;
      RECT 284.9 0.52 285.16 13.45 ;
      RECT 285.375 384.61 285.575 385.34 ;
      RECT 285.92 0.155 286.69 0.445 ;
      RECT 285.92 0.155 286.18 8.665 ;
      RECT 286.43 0.155 286.69 8.665 ;
      RECT 285.41 0.52 285.67 11.315 ;
      RECT 285.785 384.61 286.145 385.34 ;
      RECT 286.355 384.61 286.555 385.34 ;
      RECT 286.94 0.52 287.2 9.955 ;
      RECT 287.01 384.61 287.21 385.34 ;
      RECT 287.42 384.61 287.78 385.34 ;
      RECT 288.075 384.61 288.275 385.34 ;
      RECT 288.57 384.61 288.93 385.34 ;
      RECT 288.98 0.3 289.24 8.7 ;
      RECT 289.14 384.61 289.34 385.34 ;
      RECT 289.795 384.61 289.995 385.34 ;
      RECT 289.49 0.18 290.26 0.88 ;
      RECT 290.205 384.61 290.565 385.34 ;
      RECT 290.775 384.61 290.975 385.34 ;
      RECT 291.43 384.61 291.63 385.34 ;
      RECT 291.685 0.52 291.945 6.28 ;
      RECT 291.84 384.61 292.2 385.34 ;
      RECT 292.495 384.61 292.695 385.34 ;
      RECT 293.06 0.52 293.32 5.57 ;
      RECT 292.99 384.61 293.35 385.34 ;
      RECT 293.56 384.61 293.76 385.34 ;
      RECT 293.57 0.3 293.83 5.235 ;
      RECT 294.08 0.52 294.34 7.78 ;
      RECT 294.215 384.61 294.415 385.34 ;
      RECT 294.625 384.61 294.985 385.34 ;
      RECT 294.93 0.52 295.19 4.315 ;
      RECT 295.195 384.61 295.395 385.34 ;
      RECT 295.85 384.61 296.05 385.34 ;
      RECT 296.105 0.52 296.365 2.82 ;
      RECT 296.26 384.61 296.62 385.34 ;
      RECT 296.915 384.61 297.115 385.34 ;
      RECT 297.41 384.61 297.77 385.34 ;
      RECT 298.345 0.18 299.115 0.88 ;
      RECT 298.345 0.18 298.605 12.9 ;
      RECT 298.855 0.18 299.115 12.9 ;
      RECT 297.635 0.52 297.895 2.82 ;
      RECT 297.98 384.61 298.18 385.34 ;
      RECT 299.365 0.155 300.135 0.445 ;
      RECT 299.365 0.155 299.625 13.21 ;
      RECT 299.875 0.155 300.135 13.21 ;
      RECT 298.635 384.61 298.835 385.34 ;
      RECT 299.045 384.61 299.405 385.34 ;
      RECT 299.615 384.61 299.815 385.34 ;
      RECT 300.27 384.61 300.47 385.34 ;
      RECT 300.68 384.61 301.04 385.34 ;
      RECT 301.335 384.61 301.535 385.34 ;
      RECT 301.83 384.61 302.19 385.34 ;
      RECT 302.07 0.52 302.33 14.115 ;
      RECT 302.4 384.61 302.6 385.34 ;
      RECT 302.58 0.52 302.84 13.45 ;
      RECT 303.055 384.61 303.255 385.34 ;
      RECT 303.6 0.155 304.37 0.445 ;
      RECT 303.6 0.155 303.86 8.665 ;
      RECT 304.11 0.155 304.37 8.665 ;
      RECT 303.09 0.52 303.35 11.315 ;
      RECT 303.465 384.61 303.825 385.34 ;
      RECT 304.035 384.61 304.235 385.34 ;
      RECT 304.62 0.52 304.88 9.955 ;
      RECT 304.69 384.61 304.89 385.34 ;
      RECT 305.1 384.61 305.46 385.34 ;
      RECT 305.755 384.61 305.955 385.34 ;
      RECT 306.25 384.61 306.61 385.34 ;
      RECT 306.66 0.3 306.92 8.7 ;
      RECT 306.82 384.61 307.02 385.34 ;
      RECT 307.475 384.61 307.675 385.34 ;
      RECT 307.17 0.18 307.94 0.88 ;
      RECT 307.885 384.61 308.245 385.34 ;
      RECT 308.455 384.61 308.655 385.34 ;
      RECT 309.11 384.61 309.31 385.34 ;
      RECT 309.365 0.52 309.625 6.28 ;
      RECT 309.52 384.61 309.88 385.34 ;
      RECT 310.175 384.61 310.375 385.34 ;
      RECT 310.74 0.52 311 5.57 ;
      RECT 310.67 384.61 311.03 385.34 ;
      RECT 311.24 384.61 311.44 385.34 ;
      RECT 311.25 0.3 311.51 5.235 ;
      RECT 311.76 0.52 312.02 7.78 ;
      RECT 311.895 384.61 312.095 385.34 ;
      RECT 312.305 384.61 312.665 385.34 ;
      RECT 312.61 0.52 312.87 4.315 ;
      RECT 312.875 384.61 313.075 385.34 ;
      RECT 313.53 384.61 313.73 385.34 ;
      RECT 313.785 0.52 314.045 2.82 ;
      RECT 313.94 384.61 314.3 385.34 ;
      RECT 314.595 384.61 314.795 385.34 ;
      RECT 315.09 384.61 315.45 385.34 ;
      RECT 316.025 0.18 316.795 0.88 ;
      RECT 316.025 0.18 316.285 12.9 ;
      RECT 316.535 0.18 316.795 12.9 ;
      RECT 315.315 0.52 315.575 2.82 ;
      RECT 315.66 384.61 315.86 385.34 ;
      RECT 317.045 0.155 317.815 0.445 ;
      RECT 317.045 0.155 317.305 13.21 ;
      RECT 317.555 0.155 317.815 13.21 ;
      RECT 316.315 384.61 316.515 385.34 ;
      RECT 316.725 384.61 317.085 385.34 ;
      RECT 317.295 384.61 317.495 385.34 ;
      RECT 317.95 384.61 318.15 385.34 ;
      RECT 318.36 384.61 318.72 385.34 ;
      RECT 319.015 384.61 319.215 385.34 ;
      RECT 319.51 384.61 319.87 385.34 ;
      RECT 319.75 0.52 320.01 14.115 ;
      RECT 320.08 384.61 320.28 385.34 ;
      RECT 320.26 0.52 320.52 13.45 ;
      RECT 320.735 384.61 320.935 385.34 ;
      RECT 321.28 0.155 322.05 0.445 ;
      RECT 321.28 0.155 321.54 8.665 ;
      RECT 321.79 0.155 322.05 8.665 ;
      RECT 320.77 0.52 321.03 11.315 ;
      RECT 321.145 384.61 321.505 385.34 ;
      RECT 321.715 384.61 321.915 385.34 ;
      RECT 322.3 0.52 322.56 9.955 ;
      RECT 322.37 384.61 322.57 385.34 ;
      RECT 322.78 384.61 323.14 385.34 ;
      RECT 323.435 384.61 323.635 385.34 ;
      RECT 323.93 384.61 324.29 385.34 ;
      RECT 324.34 0.3 324.6 8.7 ;
      RECT 324.5 384.61 324.7 385.34 ;
      RECT 325.155 384.61 325.355 385.34 ;
      RECT 324.85 0.18 325.62 0.88 ;
      RECT 325.565 384.61 325.925 385.34 ;
      RECT 326.135 384.61 326.335 385.34 ;
      RECT 326.79 384.61 326.99 385.34 ;
      RECT 327.045 0.52 327.305 6.28 ;
      RECT 327.2 384.61 327.56 385.34 ;
      RECT 327.855 384.61 328.055 385.34 ;
      RECT 328.42 0.52 328.68 5.57 ;
      RECT 328.35 384.61 328.71 385.34 ;
      RECT 328.92 384.61 329.12 385.34 ;
      RECT 328.93 0.3 329.19 5.235 ;
      RECT 329.44 0.52 329.7 7.78 ;
      RECT 329.575 384.61 329.775 385.34 ;
      RECT 329.985 384.61 330.345 385.34 ;
      RECT 330.29 0.52 330.55 4.315 ;
      RECT 330.555 384.61 330.755 385.34 ;
      RECT 331.21 384.61 331.41 385.34 ;
      RECT 331.465 0.52 331.725 2.82 ;
      RECT 331.62 384.61 331.98 385.34 ;
      RECT 332.275 384.61 332.475 385.34 ;
      RECT 332.77 384.61 333.13 385.34 ;
      RECT 333.705 0.18 334.475 0.88 ;
      RECT 333.705 0.18 333.965 12.9 ;
      RECT 334.215 0.18 334.475 12.9 ;
      RECT 332.995 0.52 333.255 2.82 ;
      RECT 333.34 384.61 333.54 385.34 ;
      RECT 334.725 0.155 335.495 0.445 ;
      RECT 334.725 0.155 334.985 13.21 ;
      RECT 335.235 0.155 335.495 13.21 ;
      RECT 333.995 384.61 334.195 385.34 ;
      RECT 334.405 384.61 334.765 385.34 ;
      RECT 334.975 384.61 335.175 385.34 ;
      RECT 335.63 384.61 335.83 385.34 ;
      RECT 336.04 384.61 336.4 385.34 ;
      RECT 336.695 384.61 336.895 385.34 ;
      RECT 337.19 384.61 337.55 385.34 ;
      RECT 337.43 0.52 337.69 14.115 ;
      RECT 337.76 384.61 337.96 385.34 ;
      RECT 337.94 0.52 338.2 13.45 ;
      RECT 338.415 384.61 338.615 385.34 ;
      RECT 338.96 0.155 339.73 0.445 ;
      RECT 338.96 0.155 339.22 8.665 ;
      RECT 339.47 0.155 339.73 8.665 ;
      RECT 338.45 0.52 338.71 11.315 ;
      RECT 338.825 384.61 339.185 385.34 ;
      RECT 339.395 384.61 339.595 385.34 ;
      RECT 339.98 0.52 340.24 9.955 ;
      RECT 340.05 384.61 340.25 385.34 ;
      RECT 340.46 384.61 340.82 385.34 ;
      RECT 341.115 384.61 341.315 385.34 ;
      RECT 341.61 384.61 341.97 385.34 ;
      RECT 342.02 0.3 342.28 8.7 ;
      RECT 342.18 384.61 342.38 385.34 ;
      RECT 342.835 384.61 343.035 385.34 ;
      RECT 342.53 0.18 343.3 0.88 ;
      RECT 343.245 384.61 343.605 385.34 ;
      RECT 343.815 384.61 344.015 385.34 ;
      RECT 344.47 384.61 344.67 385.34 ;
      RECT 344.725 0.52 344.985 6.28 ;
      RECT 344.88 384.61 345.24 385.34 ;
      RECT 345.535 384.61 345.735 385.34 ;
      RECT 346.1 0.52 346.36 5.57 ;
      RECT 346.03 384.61 346.39 385.34 ;
      RECT 346.6 384.61 346.8 385.34 ;
      RECT 346.61 0.3 346.87 5.235 ;
      RECT 347.12 0.52 347.38 7.78 ;
      RECT 347.255 384.61 347.455 385.34 ;
      RECT 347.665 384.61 348.025 385.34 ;
      RECT 347.97 0.52 348.23 4.315 ;
      RECT 348.235 384.61 348.435 385.34 ;
      RECT 348.89 384.61 349.09 385.34 ;
      RECT 349.145 0.52 349.405 2.82 ;
      RECT 349.3 384.61 349.66 385.34 ;
      RECT 349.955 384.61 350.155 385.34 ;
      RECT 350.45 384.61 350.81 385.34 ;
      RECT 351.385 0.18 352.155 0.88 ;
      RECT 351.385 0.18 351.645 12.9 ;
      RECT 351.895 0.18 352.155 12.9 ;
      RECT 350.675 0.52 350.935 2.82 ;
      RECT 351.02 384.61 351.22 385.34 ;
      RECT 352.405 0.155 353.175 0.445 ;
      RECT 352.405 0.155 352.665 13.21 ;
      RECT 352.915 0.155 353.175 13.21 ;
      RECT 351.675 384.61 351.875 385.34 ;
      RECT 352.085 384.61 352.445 385.34 ;
      RECT 352.655 384.61 352.855 385.34 ;
      RECT 353.31 384.61 353.51 385.34 ;
      RECT 353.72 384.61 354.08 385.34 ;
      RECT 354.375 384.61 354.575 385.34 ;
      RECT 354.87 384.61 355.23 385.34 ;
      RECT 355.11 0.52 355.37 14.115 ;
      RECT 355.44 384.61 355.64 385.34 ;
      RECT 355.62 0.52 355.88 13.45 ;
      RECT 356.095 384.61 356.295 385.34 ;
      RECT 356.64 0.155 357.41 0.445 ;
      RECT 356.64 0.155 356.9 8.665 ;
      RECT 357.15 0.155 357.41 8.665 ;
      RECT 356.13 0.52 356.39 11.315 ;
      RECT 356.505 384.61 356.865 385.34 ;
      RECT 357.075 384.61 357.275 385.34 ;
      RECT 357.66 0.52 357.92 9.955 ;
      RECT 357.73 384.61 357.93 385.34 ;
      RECT 358.14 384.61 358.5 385.34 ;
      RECT 358.795 384.61 358.995 385.34 ;
      RECT 359.29 384.61 359.65 385.34 ;
      RECT 359.7 0.3 359.96 8.7 ;
      RECT 359.86 384.61 360.06 385.34 ;
      RECT 360.515 384.61 360.715 385.34 ;
      RECT 360.21 0.18 360.98 0.88 ;
      RECT 360.925 384.61 361.285 385.34 ;
      RECT 361.495 384.61 361.695 385.34 ;
      RECT 362.15 384.61 362.35 385.34 ;
      RECT 362.405 0.52 362.665 6.28 ;
      RECT 362.56 384.61 362.92 385.34 ;
      RECT 363.215 384.61 363.415 385.34 ;
      RECT 363.78 0.52 364.04 5.57 ;
      RECT 363.71 384.61 364.07 385.34 ;
      RECT 364.28 384.61 364.48 385.34 ;
      RECT 364.29 0.3 364.55 5.235 ;
      RECT 364.8 0.52 365.06 7.78 ;
      RECT 364.935 384.61 365.135 385.34 ;
      RECT 365.345 384.61 365.705 385.34 ;
      RECT 365.65 0.52 365.91 4.315 ;
      RECT 365.915 384.61 366.115 385.34 ;
      RECT 366.57 384.61 366.77 385.34 ;
      RECT 366.825 0.52 367.085 2.82 ;
      RECT 366.98 384.61 367.34 385.34 ;
      RECT 367.635 384.61 367.835 385.34 ;
      RECT 368.13 384.61 368.49 385.34 ;
      RECT 369.065 0.18 369.835 0.88 ;
      RECT 369.065 0.18 369.325 12.9 ;
      RECT 369.575 0.18 369.835 12.9 ;
      RECT 368.355 0.52 368.615 2.82 ;
      RECT 368.7 384.61 368.9 385.34 ;
      RECT 370.085 0.155 370.855 0.445 ;
      RECT 370.085 0.155 370.345 13.21 ;
      RECT 370.595 0.155 370.855 13.21 ;
      RECT 369.355 384.61 369.555 385.34 ;
      RECT 369.765 384.61 370.125 385.34 ;
      RECT 370.335 384.61 370.535 385.34 ;
      RECT 370.99 384.61 371.19 385.34 ;
      RECT 371.4 384.61 371.76 385.34 ;
      RECT 372.055 384.61 372.255 385.34 ;
      RECT 372.55 384.61 372.91 385.34 ;
      RECT 372.79 0.52 373.05 14.115 ;
      RECT 373.12 384.61 373.32 385.34 ;
      RECT 373.3 0.52 373.56 13.45 ;
      RECT 373.775 384.61 373.975 385.34 ;
      RECT 374.32 0.155 375.09 0.445 ;
      RECT 374.32 0.155 374.58 8.665 ;
      RECT 374.83 0.155 375.09 8.665 ;
      RECT 373.81 0.52 374.07 11.315 ;
      RECT 374.185 384.61 374.545 385.34 ;
      RECT 374.755 384.61 374.955 385.34 ;
      RECT 375.34 0.52 375.6 9.955 ;
      RECT 375.41 384.61 375.61 385.34 ;
      RECT 375.82 384.61 376.18 385.34 ;
      RECT 376.475 384.61 376.675 385.34 ;
      RECT 376.97 384.61 377.33 385.34 ;
      RECT 377.38 0.3 377.64 8.7 ;
      RECT 377.54 384.61 377.74 385.34 ;
      RECT 378.195 384.61 378.395 385.34 ;
      RECT 377.89 0.18 378.66 0.88 ;
      RECT 378.605 384.61 378.965 385.34 ;
      RECT 379.175 384.61 379.375 385.34 ;
      RECT 379.83 384.61 380.03 385.34 ;
      RECT 380.085 0.52 380.345 6.28 ;
      RECT 380.24 384.61 380.6 385.34 ;
      RECT 380.895 384.61 381.095 385.34 ;
      RECT 381.46 0.52 381.72 5.57 ;
      RECT 381.39 384.61 381.75 385.34 ;
      RECT 381.96 384.61 382.16 385.34 ;
      RECT 381.97 0.3 382.23 5.235 ;
      RECT 382.48 0.52 382.74 7.78 ;
      RECT 382.615 384.61 382.815 385.34 ;
      RECT 383.025 384.61 383.385 385.34 ;
      RECT 383.33 0.52 383.59 4.315 ;
      RECT 383.595 384.61 383.795 385.34 ;
      RECT 384.25 384.61 384.45 385.34 ;
      RECT 384.505 0.52 384.765 2.82 ;
      RECT 384.66 384.61 385.02 385.34 ;
      RECT 385.315 384.61 385.515 385.34 ;
      RECT 385.81 384.61 386.17 385.34 ;
      RECT 386.745 0.18 387.515 0.88 ;
      RECT 386.745 0.18 387.005 12.9 ;
      RECT 387.255 0.18 387.515 12.9 ;
      RECT 386.035 0.52 386.295 2.82 ;
      RECT 386.38 384.61 386.58 385.34 ;
      RECT 387.765 0.155 388.535 0.445 ;
      RECT 387.765 0.155 388.025 13.21 ;
      RECT 388.275 0.155 388.535 13.21 ;
      RECT 387.035 384.61 387.235 385.34 ;
      RECT 387.445 384.61 387.805 385.34 ;
      RECT 388.015 384.61 388.215 385.34 ;
      RECT 388.67 384.61 388.87 385.34 ;
      RECT 389.08 384.61 389.44 385.34 ;
      RECT 389.735 384.61 389.935 385.34 ;
      RECT 390.23 384.61 390.59 385.34 ;
      RECT 390.47 0.52 390.73 14.115 ;
      RECT 390.8 384.61 391 385.34 ;
      RECT 390.98 0.52 391.24 13.45 ;
      RECT 391.455 384.61 391.655 385.34 ;
      RECT 392 0.155 392.77 0.445 ;
      RECT 392 0.155 392.26 8.665 ;
      RECT 392.51 0.155 392.77 8.665 ;
      RECT 391.49 0.52 391.75 11.315 ;
      RECT 391.865 384.61 392.225 385.34 ;
      RECT 392.435 384.61 392.635 385.34 ;
      RECT 393.02 0.52 393.28 9.955 ;
      RECT 393.09 384.61 393.29 385.34 ;
      RECT 393.5 384.61 393.86 385.34 ;
      RECT 394.155 384.61 394.355 385.34 ;
      RECT 394.65 384.61 395.01 385.34 ;
      RECT 395.06 0.3 395.32 8.7 ;
      RECT 395.22 384.61 395.42 385.34 ;
      RECT 395.875 384.61 396.075 385.34 ;
      RECT 395.57 0.18 396.34 0.88 ;
      RECT 396.285 384.61 396.645 385.34 ;
      RECT 396.855 384.61 397.055 385.34 ;
      RECT 397.51 384.61 397.71 385.34 ;
      RECT 397.765 0.52 398.025 6.28 ;
      RECT 397.92 384.61 398.28 385.34 ;
      RECT 398.575 384.61 398.775 385.34 ;
      RECT 399.14 0.52 399.4 5.57 ;
      RECT 399.07 384.61 399.43 385.34 ;
      RECT 399.64 384.61 399.84 385.34 ;
      RECT 399.65 0.3 399.91 5.235 ;
      RECT 400.16 0.52 400.42 7.78 ;
      RECT 400.295 384.61 400.495 385.34 ;
      RECT 400.705 384.61 401.065 385.34 ;
      RECT 401.275 384.61 401.475 385.34 ;
      RECT 402.1 53.41 402.3 385.34 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 398.285 0 398.88 385.37 ;
      RECT 399.65 0.3 399.91 385.37 ;
      RECT 400.68 0 402.61 385.37 ;
      RECT 0 0.52 402.61 385.37 ;
      RECT 393.54 0 397.505 385.37 ;
      RECT 392 0.155 392.77 385.37 ;
      RECT 386.555 0 390.21 385.37 ;
      RECT 385.025 0 385.775 385.37 ;
      RECT 383.85 0 384.245 385.37 ;
      RECT 381.97 0.3 382.23 385.37 ;
      RECT 380.605 0 381.2 385.37 ;
      RECT 375.86 0 379.825 385.37 ;
      RECT 374.32 0.155 375.09 385.37 ;
      RECT 368.875 0 372.53 385.37 ;
      RECT 367.345 0 368.095 385.37 ;
      RECT 366.17 0 366.565 385.37 ;
      RECT 364.29 0.3 364.55 385.37 ;
      RECT 362.925 0 363.52 385.37 ;
      RECT 358.18 0 362.145 385.37 ;
      RECT 356.64 0.155 357.41 385.37 ;
      RECT 351.195 0 354.85 385.37 ;
      RECT 349.665 0 350.415 385.37 ;
      RECT 348.49 0 348.885 385.37 ;
      RECT 346.61 0.3 346.87 385.37 ;
      RECT 345.245 0 345.84 385.37 ;
      RECT 340.5 0 344.465 385.37 ;
      RECT 338.96 0.155 339.73 385.37 ;
      RECT 333.515 0 337.17 385.37 ;
      RECT 331.985 0 332.735 385.37 ;
      RECT 330.81 0 331.205 385.37 ;
      RECT 328.93 0.3 329.19 385.37 ;
      RECT 327.565 0 328.16 385.37 ;
      RECT 322.82 0 326.785 385.37 ;
      RECT 321.28 0.155 322.05 385.37 ;
      RECT 315.835 0 319.49 385.37 ;
      RECT 314.305 0 315.055 385.37 ;
      RECT 313.13 0 313.525 385.37 ;
      RECT 311.25 0.3 311.51 385.37 ;
      RECT 309.885 0 310.48 385.37 ;
      RECT 305.14 0 309.105 385.37 ;
      RECT 303.6 0.155 304.37 385.37 ;
      RECT 298.155 0 301.81 385.37 ;
      RECT 296.625 0 297.375 385.37 ;
      RECT 295.45 0 295.845 385.37 ;
      RECT 293.57 0.3 293.83 385.37 ;
      RECT 292.205 0 292.8 385.37 ;
      RECT 287.46 0 291.425 385.37 ;
      RECT 285.92 0.155 286.69 385.37 ;
      RECT 280.475 0 284.13 385.37 ;
      RECT 278.945 0 279.695 385.37 ;
      RECT 277.77 0 278.165 385.37 ;
      RECT 275.89 0.3 276.15 385.37 ;
      RECT 274.525 0 275.12 385.37 ;
      RECT 269.78 0 273.745 385.37 ;
      RECT 268.24 0.155 269.01 385.37 ;
      RECT 262.795 0 266.45 385.37 ;
      RECT 261.265 0 262.015 385.37 ;
      RECT 260.09 0 260.485 385.37 ;
      RECT 237.285 0.18 259.31 385.37 ;
      RECT 237.295 0 259.31 385.37 ;
      RECT 232.695 0.3 236.525 385.37 ;
      RECT 230.655 0.18 231.425 385.37 ;
      RECT 224.025 0.3 225.305 385.37 ;
      RECT 221.475 0.3 222.755 385.37 ;
      RECT 219.945 0.3 220.205 385.37 ;
      RECT 216.885 0.3 217.145 385.37 ;
      RECT 215.355 0.3 215.615 385.37 ;
      RECT 207.195 0.3 214.085 385.37 ;
      RECT 197.705 0 204.905 385.37 ;
      RECT 188.525 0.3 195.415 385.37 ;
      RECT 188.535 0 195.415 385.37 ;
      RECT 186.995 0.3 187.255 385.37 ;
      RECT 185.465 0.3 185.725 385.37 ;
      RECT 182.405 0.3 182.665 385.37 ;
      RECT 179.855 0.3 181.135 385.37 ;
      RECT 177.305 0.3 178.585 385.37 ;
      RECT 171.185 0.18 171.955 385.37 ;
      RECT 166.085 0.3 169.915 385.37 ;
      RECT 143.3 0.18 165.325 385.37 ;
      RECT 142.125 0 142.52 385.37 ;
      RECT 140.595 0 141.345 385.37 ;
      RECT 136.16 0 139.815 385.37 ;
      RECT 133.6 0.155 134.37 385.37 ;
      RECT 128.865 0 132.83 385.37 ;
      RECT 127.49 0 128.085 385.37 ;
      RECT 126.46 0.3 126.72 385.37 ;
      RECT 124.445 0 124.84 385.37 ;
      RECT 122.915 0 123.665 385.37 ;
      RECT 118.48 0 122.135 385.37 ;
      RECT 115.92 0.155 116.69 385.37 ;
      RECT 111.185 0 115.15 385.37 ;
      RECT 109.81 0 110.405 385.37 ;
      RECT 108.78 0.3 109.04 385.37 ;
      RECT 106.765 0 107.16 385.37 ;
      RECT 105.235 0 105.985 385.37 ;
      RECT 100.8 0 104.455 385.37 ;
      RECT 98.24 0.155 99.01 385.37 ;
      RECT 93.505 0 97.47 385.37 ;
      RECT 92.13 0 92.725 385.37 ;
      RECT 91.1 0.3 91.36 385.37 ;
      RECT 89.085 0 89.48 385.37 ;
      RECT 87.555 0 88.305 385.37 ;
      RECT 83.12 0 86.775 385.37 ;
      RECT 80.56 0.155 81.33 385.37 ;
      RECT 75.825 0 79.79 385.37 ;
      RECT 74.45 0 75.045 385.37 ;
      RECT 73.42 0.3 73.68 385.37 ;
      RECT 71.405 0 71.8 385.37 ;
      RECT 69.875 0 70.625 385.37 ;
      RECT 65.44 0 69.095 385.37 ;
      RECT 62.88 0.155 63.65 385.37 ;
      RECT 58.145 0 62.11 385.37 ;
      RECT 56.77 0 57.365 385.37 ;
      RECT 55.74 0.3 56 385.37 ;
      RECT 53.725 0 54.12 385.37 ;
      RECT 52.195 0 52.945 385.37 ;
      RECT 47.76 0 51.415 385.37 ;
      RECT 45.2 0.155 45.97 385.37 ;
      RECT 40.465 0 44.43 385.37 ;
      RECT 39.09 0 39.685 385.37 ;
      RECT 38.06 0.3 38.32 385.37 ;
      RECT 36.045 0 36.44 385.37 ;
      RECT 34.515 0 35.265 385.37 ;
      RECT 30.08 0 33.735 385.37 ;
      RECT 27.52 0.155 28.29 385.37 ;
      RECT 22.785 0 26.75 385.37 ;
      RECT 21.41 0 22.005 385.37 ;
      RECT 20.38 0.3 20.64 385.37 ;
      RECT 18.365 0 18.76 385.37 ;
      RECT 16.835 0 17.585 385.37 ;
      RECT 12.4 0 16.055 385.37 ;
      RECT 9.84 0.155 10.61 385.37 ;
      RECT 5.105 0 9.07 385.37 ;
      RECT 3.73 0 4.325 385.37 ;
      RECT 2.7 0.3 2.96 385.37 ;
      RECT 0 0 1.93 385.37 ;
      RECT 399.66 0 399.9 385.37 ;
      RECT 381.98 0 382.22 385.37 ;
      RECT 364.3 0 364.54 385.37 ;
      RECT 346.62 0 346.86 385.37 ;
      RECT 328.94 0 329.18 385.37 ;
      RECT 311.26 0 311.5 385.37 ;
      RECT 293.58 0 293.82 385.37 ;
      RECT 275.9 0 276.14 385.37 ;
      RECT 232.705 0 236.515 385.37 ;
      RECT 224.035 0 225.295 385.37 ;
      RECT 221.485 0 222.745 385.37 ;
      RECT 219.955 0 220.195 385.37 ;
      RECT 216.895 0 217.135 385.37 ;
      RECT 215.365 0 215.605 385.37 ;
      RECT 207.195 0 214.075 385.37 ;
      RECT 187.005 0 187.245 385.37 ;
      RECT 185.475 0 185.715 385.37 ;
      RECT 182.415 0 182.655 385.37 ;
      RECT 179.865 0 181.125 385.37 ;
      RECT 177.315 0 178.575 385.37 ;
      RECT 166.095 0 169.905 385.37 ;
      RECT 126.47 0 126.71 385.37 ;
      RECT 108.79 0 109.03 385.37 ;
      RECT 91.11 0 91.35 385.37 ;
      RECT 73.43 0 73.67 385.37 ;
      RECT 55.75 0 55.99 385.37 ;
      RECT 38.07 0 38.31 385.37 ;
      RECT 20.39 0 20.63 385.37 ;
      RECT 2.71 0 2.95 385.37 ;
      RECT 230.665 0 231.415 385.37 ;
      RECT 171.195 0 171.945 385.37 ;
      RECT 143.3 0 165.315 385.37 ;
      RECT 392.01 0 392.76 385.37 ;
      RECT 374.33 0 375.08 385.37 ;
      RECT 356.65 0 357.4 385.37 ;
      RECT 338.97 0 339.72 385.37 ;
      RECT 321.29 0 322.04 385.37 ;
      RECT 303.61 0 304.36 385.37 ;
      RECT 285.93 0 286.68 385.37 ;
      RECT 268.25 0 269 385.37 ;
      RECT 133.61 0 134.36 385.37 ;
      RECT 115.93 0 116.68 385.37 ;
      RECT 98.25 0 99 385.37 ;
      RECT 80.57 0 81.32 385.37 ;
      RECT 62.89 0 63.64 385.37 ;
      RECT 45.21 0 45.96 385.37 ;
      RECT 27.53 0 28.28 385.37 ;
      RECT 9.85 0 10.6 385.37 ;
    LAYER Metal3 ;
      RECT 0 0 402.61 385.37 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 241.595 0 259.185 385.37 ;
      RECT 236.445 0 238.265 385.37 ;
      RECT 231.295 0 233.115 385.37 ;
      RECT 396.725 0 402.61 385.37 ;
      RECT 387.885 0 391.785 385.37 ;
      RECT 387.885 47.305 402.61 53.15 ;
      RECT 379.045 0 382.945 385.37 ;
      RECT 370.205 0 374.105 385.37 ;
      RECT 370.205 47.305 382.945 53.15 ;
      RECT 361.365 0 365.265 385.37 ;
      RECT 352.525 0 356.425 385.37 ;
      RECT 352.525 47.305 365.265 53.15 ;
      RECT 343.685 0 347.585 385.37 ;
      RECT 334.845 0 338.745 385.37 ;
      RECT 334.845 47.305 347.585 53.15 ;
      RECT 326.005 0 329.905 385.37 ;
      RECT 317.165 0 321.065 385.37 ;
      RECT 317.165 47.305 329.905 53.15 ;
      RECT 308.325 0 312.225 385.37 ;
      RECT 299.485 0 303.385 385.37 ;
      RECT 299.485 47.305 312.225 53.15 ;
      RECT 290.645 0 294.545 385.37 ;
      RECT 281.805 0 285.705 385.37 ;
      RECT 281.805 47.305 294.545 53.15 ;
      RECT 272.965 0 276.865 385.37 ;
      RECT 264.125 0 268.025 385.37 ;
      RECT 264.125 47.305 276.865 53.15 ;
      RECT 226.145 0 227.965 385.37 ;
      RECT 220.995 0 222.815 385.37 ;
      RECT 215.845 0 217.665 385.37 ;
      RECT 210.695 0 212.515 385.37 ;
      RECT 205.545 0 207.365 385.37 ;
      RECT 200.395 0 202.215 385.37 ;
      RECT 195.245 0 197.065 385.37 ;
      RECT 190.095 0 191.915 385.37 ;
      RECT 184.945 0 186.765 385.37 ;
      RECT 179.795 0 181.615 385.37 ;
      RECT 174.645 0 176.465 385.37 ;
      RECT 169.495 0 171.315 385.37 ;
      RECT 164.345 0 166.165 385.37 ;
      RECT 143.425 0 161.015 385.37 ;
      RECT 134.585 0 138.485 385.37 ;
      RECT 125.745 0 129.645 385.37 ;
      RECT 125.745 47.305 138.485 53.15 ;
      RECT 116.905 0 120.805 385.37 ;
      RECT 108.065 0 111.965 385.37 ;
      RECT 108.065 47.305 120.805 53.15 ;
      RECT 99.225 0 103.125 385.37 ;
      RECT 90.385 0 94.285 385.37 ;
      RECT 90.385 47.305 103.125 53.15 ;
      RECT 81.545 0 85.445 385.37 ;
      RECT 72.705 0 76.605 385.37 ;
      RECT 72.705 47.305 85.445 53.15 ;
      RECT 63.865 0 67.765 385.37 ;
      RECT 55.025 0 58.925 385.37 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 385.37 ;
      RECT 37.345 0 41.245 385.37 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 385.37 ;
      RECT 19.665 0 23.565 385.37 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 385.37 ;
      RECT 0 0 5.885 385.37 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_1024x16_c2_bm_bist

END LIBRARY
