* ------------------------------------------------------
*
*		Copyright 2025 IHP PDK Authors
*
*		Licensed under the Apache License, Version 2.0 (the "License");
*		you may not use this file except in compliance with the License.
*		You may obtain a copy of the License at
*		
*		   https://www.apache.org/licenses/LICENSE-2.0
*		
*		Unless required by applicable law or agreed to in writing, software
*		distributed under the License is distributed on an "AS IS" BASIS,
*		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*		See the License for the specific language governing permissions and
*		limitations under the License.
*		
*		Generated on Wed Aug 27 13:36:37 2025		
*
* ------------------------------------------------------ 

.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR LWL NW PW VDD VSS
MN1 VSS LWL VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS net9 VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<14> A_WL<14> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<13> A_WL<13> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<12> A_WL<12> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<11> A_WL<11> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<10> A_WL<10> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<9> A_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<8> A_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<7> A_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<6> A_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<5> A_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<4> A_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<3> A_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<2> A_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<1> A_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
XI0<0> A_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_CELL BLC_BOT BLC_TOP BLT_BOT BLT_TOP LWL NW PW 
+ RWL VDD VSS
MN0 NC NT VSS PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN1 NT NC VSS PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN3 NC RWL BLC_TOP PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 BLT_BOT LWL NT PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW sg13_lv_pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW sg13_lv_pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R1 BLC_BOT BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 BLT_BOT BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 RWL LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE 
+ VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_RWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_RWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_RWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_RWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_RWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_RWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_RWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_RWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_RWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_RWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_RWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_RWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_RWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_RWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_RWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_RWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX4 A Z VDD VSS
MN0 net9 A VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 Z net9 VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 net9 A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net9 VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX4 A Z VDD VSS
MN1 Z net6 VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net6 A VSS VSS sg13_lv_nmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net6 VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 A VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP8 VDD VSS
MN0 vss_r vdd_r VSS VSS sg13_lv_nmos m=1 w=4.98u l=130.00n ng=6 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD sg13_lv_pmos m=1 w=6.48u l=385.000n ng=4 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_LHPQX2 CP D Q VDD VSS
MN3 QIN CPN net14 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net14 net10 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN5 net21 D VSS VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 QIN CP net21 VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net10 QIN VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 Q QIN VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 QIN CP net16 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 CPN CP VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 Q QIN VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 net10 QIN VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net16 net10 VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 QIN CPN net20 VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP5 net20 D VDD VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND2X2 A B Z VDD VSS
MP1 Z B VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B net7 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net7 A VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4 A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX2 A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX2 A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND3X2 A B C Z VDD VSS
MP2 Z A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z B VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z C VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 net12 B net16 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C net12 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net16 A VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NOR3X2 A B C Z VDD VSS
MP0 net13 A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 Z C net10 VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 net10 B net13 VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 Z B VSS VSS sg13_lv_nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C VSS VSS sg13_lv_nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN2 Z A VSS VSS sg13_lv_nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP4 VDD VSS
MN0 vss_r vdd_r VSS VSS sg13_lv_nmos m=1 w=2.49u l=130.00n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD sg13_lv_pmos m=1 w=3.24u l=385.000n ng=2 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET2RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
.ENDS
.SUBCKT RSC_IHPSG13_CINVX8 A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_DFNQMX2IX1 BE BI CN D QI QIN VDD VSS
MN15 net026 BI VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN14 MXI_OUT BE net026 VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net025 D VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 MXI_OUT BEN net025 VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QI CNN net21 VSS sg13_lv_nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 nrs=0
MN11 net21 QI_MS VSS VSS sg13_lv_nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS sg13_lv_nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 MXI_OUT VSS VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN_MS CN net37 VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QI CN net25 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN4 net25 QIN VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 QIN QI VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN13 BEN BE VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP15 MXI_OUT BEN net027 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP14 net027 BI VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP1 MXI_OUT BE net024 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net024 D VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP13 BEN BE VDD VDD sg13_lv_pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QI CNN net27 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 net27 QIN VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP10 net36 MXI_OUT VDD VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP11 QIN_MS CNN net36 VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QIN QI VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 CNN CN VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QI CN net19 VDD sg13_lv_pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 nrs=0
MP8 net19 QI_MS VDD VDD sg13_lv_pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1 A Z VDD VSS
MN1 net010 net032 VSS VSS sg13_lv_nmos m=1 w=300.0n l=160.00n ng=1 
+ nrd=0 nrs=0
MN2 net032 A net014 VSS sg13_lv_nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN0 Z net032 net010 VSS sg13_lv_nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN3 net014 A VSS VSS sg13_lv_nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net032 net07 VDD sg13_lv_pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP3 net011 A VDD VDD sg13_lv_pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP0 net07 net032 VDD VDD sg13_lv_pmos m=1 w=720.00n l=160.00n ng=1 
+ nrd=0 nrs=0
MP2 net032 A net011 VDD sg13_lv_pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1_DUMMY A Z VDD VSS
MN0 vss_r vdd_r VSS VSS sg13_lv_nmos m=1 w=2.49u l=300.0n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD sg13_lv_pmos m=1 w=3.24u l=640.00n ng=2 nrd=0 
+ nrs=0
R0 Z A lvsres w=2.6e-07 l=6e-07
.ENDS

.SUBCKT RSC_IHPSG13_MX2IX1 A0 A1 S ZN VDD VSS
MP4 SN S VDD VDD sg13_lv_pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 ZN SN net12 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP2 net12 A1 VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 ZN S net17 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 net17 A0 VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 ZN S net13 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net15 A0 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 ZN SN net15 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RSC_IHPSG13_DFNQX2 CN D Q VDD VSS
MN0 Q QIN_SL VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QIN_SL CNN net21 VSS sg13_lv_nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN11 net21 QI_MS VSS VSS sg13_lv_nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS sg13_lv_nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 D VSS VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN8 QIN_MS CN net37 VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QIN_SL CN net25 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net25 QI_SL VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN2 QI_SL QIN_SL VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 Q QIN_SL VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QIN_SL CNN net27 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net27 QI_SL VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP10 net36 D VDD VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 QIN_MS CNN net36 VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QI_SL QIN_SL VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP12 CNN CN VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QIN_SL CN net19 VDD sg13_lv_pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP8 net19 QI_MS VDD VDD sg13_lv_pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CNAND2X2 A B Z VDD VSS
MN0 Z B net6 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net6 A VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z B VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CGATEPX4 CP E Q VDD VSS
MN1 net08 QIN VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net019 net08 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN3 QIN CP net019 VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN6 Q net015 VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 
+ nrs=0
MN5 net015 net08 net018 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN CPN net023 VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net023 E VSS VSS sg13_lv_nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net018 CP VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP3 net08 QIN VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 QIN CPN net017 VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net017 net08 VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 CPN CP VDD VDD sg13_lv_pmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP8 QIN CP net024 VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net024 E VDD VDD sg13_lv_pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net015 CP VDD VDD sg13_lv_pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 Q net015 VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 
+ nrs=0
MP5 net015 net08 VDD VDD sg13_lv_pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX8 A Z VDD VSS
MP0 net4 A VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net4 VDD VDD sg13_lv_pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MN1 Z net4 VSS VSS sg13_lv_nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MN0 net4 A VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX2 A Z VDD VSS
MN2 net4 A net9 VSS sg13_lv_nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MN0 Z net4 VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net9 A VSS VSS sg13_lv_nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MP2 net4 A net10 VDD sg13_lv_pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP1 net10 A VDD VDD sg13_lv_pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP0 Z net4 VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MX2X2 A0 A1 S Z VDD VSS
MP6 Z net010 VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 SN S VDD VDD sg13_lv_pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 net010 SN net12 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net12 A1 VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net010 S net17 VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net17 A0 VDD VDD sg13_lv_pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 Z net010 VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net010 S net13 VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net15 A0 VSS VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net010 SN net15 VSS sg13_lv_nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_AND2X2 A B Z VDD VSS
MN3 Z net6 VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net9 B VSS VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net6 B VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_TIEL Z VDD VSS
MN0 Z net2 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net2 net2 VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_XOR2X2 A B Z VDD VSS
MP8 net012 B net7 VDD sg13_lv_pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net011 net3 net012 VDD sg13_lv_pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 Z net012 VDD VDD sg13_lv_pmos m=1 w=1.535u l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net7 A VDD VDD sg13_lv_pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net011 net7 VDD VDD sg13_lv_pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 net3 B VDD VDD sg13_lv_pmos m=1 w=580.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net012 B net011 VSS sg13_lv_nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 net7 net3 net012 VSS sg13_lv_nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 Z net012 VSS VSS sg13_lv_nmos m=1 w=775.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net7 A VSS VSS sg13_lv_nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net3 B VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 net011 net7 VSS VSS sg13_lv_nmos m=1 w=555.000n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_OA12X1 A B C Z VDD VSS
MN2 net7 C VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 Z net17 VSS VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net17 B net7 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 net17 A net7 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 net24 A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 Z net17 VDD VDD sg13_lv_pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net17 B net24 VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 net17 C VDD VDD sg13_lv_pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net9 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net9 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net9 net8 VDD VSS / RSC_IHPSG13_CINVX2
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XI6 PULSE_L PULSE_H net9 VDD VSS / RSC_IHPSG13_XOR2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<3> PADR<1> PADR<0> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> PADR<1> NADR<0> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> NADR<1> PADR<0> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<1> NADR<0> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI16<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI17<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI17<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI17<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RSC_IHPSG13_NOR2X2 A B Z VDD VSS
MP1 Z B net9 VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net9 A VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 Z A VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4_WN A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BLDRV BLC BLC_SEL BLT BLT_SEL PRE_N SEL_P WR_ONE WR_ZERO 
+ VDD VSS
XCDEC SEL_P WR_ZERO BLC_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
XTDEC SEL_P WR_ONE BLT_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
MTWN BLT BLT_NMOS_DRIVE VSS VSS sg13_lv_nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWN BLC BLC_NMOS_DRIVE VSS VSS sg13_lv_nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWP BLC BLC_PMOS_DRIVE VDD VDD sg13_lv_pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTWP BLT BLT_PMOS_DRIVE VDD VDD sg13_lv_pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTSP BLT_SEL SEL_N BLT VDD sg13_lv_pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MTPR BLT PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
MCSP BLC_SEL SEL_N BLC VDD sg13_lv_pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MCPR BLC PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
XI86 SEL_P SEL_N VDD VSS / RSC_IHPSG13_INVX2
XTINV BLC_PMOS_DRIVE BLT_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
XCINV BLT_PMOS_DRIVE BLC_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RSC_IHPSG13_TIEH Z VDD VSS
MN0 net2 net2 VSS VSS sg13_lv_nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 Z net2 VDD VDD sg13_lv_pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET3RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2 CP DN DP QN QP VDD VSS
MN12 SN RN DIFFP VSS sg13_lv_nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN13 TAIL CP VSS VSS sg13_lv_nmos m=1 w=2.4u l=130.00n ng=2 nrd=0 nrs=0
MN9 DIFFP DP TAIL VSS sg13_lv_nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN10 DIFFN DN TAIL VSS sg13_lv_nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN11 RN SN DIFFN VSS sg13_lv_nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN19 net33 SN VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN20 QN QP net37 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN18 net37 RN VSS VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN17 QP QN net33 VSS sg13_lv_nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP15 SN RN VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP16 RN CP VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP14 DIFFP CP VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 RN SN VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP13 DIFFN CP VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 SN CP VDD VDD sg13_lv_pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP19 QN QP VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP20 QP SN VDD VDD sg13_lv_pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP18 QN RN VDD VDD sg13_lv_pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP17 QP QN VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX2 A Z VDD VSS
MN1 Z net4 VSS VSS sg13_lv_nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net4 A VSS VSS sg13_lv_nmos m=1 w=540.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net4 VDD VDD sg13_lv_pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net4 A VDD VDD sg13_lv_pmos m=1 w=1.1u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX4 A Z VDD VSS
MN0 Z A VSS VSS sg13_lv_nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I44 A_WCLK_B_R A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_R A_RCLK_B_L / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_R A_RCLK_L / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_R A_WCLK_B_L / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I78 A_RCLK_B_R A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_R A_RCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13_FILL4 VDD VSS
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net7<0> VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_AND2X4 A B Z VDD VSS
MN3 Z net6 VSS VSS sg13_lv_nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MN4 net9 B VSS VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 B VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DO_WRITE_P A_DI_N A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_R A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_I70<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I44 A_BM_N A_WCLK_B_R A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_ADDR_DEC<6> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_ADDR_DEC<5> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<4> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR A_WL B_WL NW PW VDD VSS
MN1 VSS A_WL VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS B_WL VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> 
+ B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> 
+ B_WL<1> B_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> B_WL<15> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<14> A_WL<14> B_WL<14> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<13> A_WL<13> B_WL<13> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<12> A_WL<12> B_WL<12> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<11> A_WL<11> B_WL<11> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<10> A_WL<10> B_WL<10> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<9> A_WL<9> B_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<8> A_WL<8> B_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<7> A_WL<7> B_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<6> A_WL<6> B_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<5> A_WL<5> B_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<4> A_WL<4> B_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<3> A_WL<3> B_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<2> A_WL<2> B_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<1> A_WL<1> B_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
XI0<0> A_WL<0> B_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_CELL A_BLC_BOT A_BLC_TOP A_BLT_BOT A_BLT_TOP 
+ A_LWL A_RWL B_BLC_BOT B_BLC_TOP B_BLT_BOT B_BLT_TOP B_LWL B_RWL NW PW VDD VSS
MN5 NC B_RWL B_BLC_BOT PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN4 B_BLT_BOT B_LWL NT PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 NC NT VSS PW sg13_lv_nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN1 NT NC VSS PW sg13_lv_nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN3 NC A_RWL A_BLC_TOP PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 A_BLT_TOP A_LWL NT PW sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW sg13_lv_pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW sg13_lv_pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R5 B_RWL B_LWL lvsres w=2.6e-07 l=6e-07
R4 B_BLC_BOT B_BLC_TOP lvsres w=2.6e-07 l=6e-07
R3 B_BLT_BOT B_BLT_TOP lvsres w=2.6e-07 l=6e-07
R1 A_BLC_BOT A_BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 A_BLT_BOT A_BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 A_RWL A_LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> B_BLC_BOT<1> 
+ B_BLC_BOT<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT_BOT<1> B_BLT_BOT<0> 
+ B_BLT_TOP<1> B_BLT_TOP<0> B_LWL<15> B_LWL<14> B_LWL<13> B_LWL<12> B_LWL<11> 
+ B_LWL<10> B_LWL<9> B_LWL<8> B_LWL<7> B_LWL<6> B_LWL<5> B_LWL<4> B_LWL<3> 
+ B_LWL<2> B_LWL<1> B_LWL<0> B_RWL<15> B_RWL<14> B_RWL<13> B_RWL<12> B_RWL<11> 
+ B_RWL<10> B_RWL<9> B_RWL<8> B_RWL<7> B_RWL<6> B_RWL<5> B_RWL<4> B_RWL<3> 
+ B_RWL<2> B_RWL<1> B_RWL<0> VDD_CORE VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_XWL<15> A_RWL<15> 
+ B_BLC_TOP<1> B_RBLC<15> B_BLT_TOP<1> B_RBLT<15> B_XWL<15> B_RWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_XWL<14> A_RWL<14> 
+ B_RBLC<14> B_RBLC<15> B_RBLT<14> B_RBLT<15> B_XWL<14> B_RWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_XWL<13> A_RWL<13> 
+ B_RBLC<14> B_RBLC<13> B_RBLT<14> B_RBLT<13> B_XWL<13> B_RWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_XWL<12> A_RWL<12> 
+ B_RBLC<12> B_RBLC<13> B_RBLT<12> B_RBLT<13> B_XWL<12> B_RWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_XWL<11> A_RWL<11> 
+ B_RBLC<12> B_RBLC<11> B_RBLT<12> B_RBLT<11> B_XWL<11> B_RWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_XWL<10> A_RWL<10> 
+ B_RBLC<10> B_RBLC<11> B_RBLT<10> B_RBLT<11> B_XWL<10> B_RWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_XWL<9> A_RWL<9> 
+ B_RBLC<10> B_RBLC<9> B_RBLT<10> B_RBLT<9> B_XWL<9> B_RWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_XWL<8> A_RWL<8> B_RBLC<8> 
+ B_RBLC<9> B_RBLT<8> B_RBLT<9> B_XWL<8> B_RWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_XWL<7> A_RWL<7> B_RBLC<8> 
+ B_RBLC<7> B_RBLT<8> B_RBLT<7> B_XWL<7> B_RWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_XWL<6> A_RWL<6> B_RBLC<6> 
+ B_RBLC<7> B_RBLT<6> B_RBLT<7> B_XWL<6> B_RWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_XWL<5> A_RWL<5> B_RBLC<6> 
+ B_RBLC<5> B_RBLT<6> B_RBLT<5> B_XWL<5> B_RWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_XWL<4> A_RWL<4> B_RBLC<4> 
+ B_RBLC<5> B_RBLT<4> B_RBLT<5> B_XWL<4> B_RWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_XWL<3> A_RWL<3> B_RBLC<4> 
+ B_RBLC<3> B_RBLT<4> B_RBLT<3> B_XWL<3> B_RWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_XWL<2> A_RWL<2> B_RBLC<2> 
+ B_RBLC<3> B_RBLT<2> B_RBLT<3> B_XWL<2> B_RWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_XWL<1> A_RWL<1> B_RBLC<2> 
+ B_RBLC<1> B_RBLT<2> B_RBLT<1> B_XWL<1> B_RWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_XWL<0> A_RWL<0> 
+ B_BLC_BOT<1> B_RBLC<1> B_BLT_BOT<1> B_RBLT<1> B_XWL<0> B_RWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> A_XWL<15> 
+ B_BLC_TOP<0> B_LBLC<15> B_BLT_TOP<0> B_LBLT<15> B_LWL<15> B_XWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> A_XWL<14> 
+ B_LBLC<14> B_LBLC<15> B_LBLT<14> B_LBLT<15> B_LWL<14> B_XWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> A_XWL<13> 
+ B_LBLC<14> B_LBLC<13> B_LBLT<14> B_LBLT<13> B_LWL<13> B_XWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> A_XWL<12> 
+ B_LBLC<12> B_LBLC<13> B_LBLT<12> B_LBLT<13> B_LWL<12> B_XWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> A_XWL<11> 
+ B_LBLC<12> B_LBLC<11> B_LBLT<12> B_LBLT<11> B_LWL<11> B_XWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> A_XWL<10> 
+ B_LBLC<10> B_LBLC<11> B_LBLT<10> B_LBLT<11> B_LWL<10> B_XWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> A_XWL<9> 
+ B_LBLC<10> B_LBLC<9> B_LBLT<10> B_LBLT<9> B_LWL<9> B_XWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> A_XWL<8> B_LBLC<8> 
+ B_LBLC<9> B_LBLT<8> B_LBLT<9> B_LWL<8> B_XWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> A_XWL<7> B_LBLC<8> 
+ B_LBLC<7> B_LBLT<8> B_LBLT<7> B_LWL<7> B_XWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> A_XWL<6> B_LBLC<6> 
+ B_LBLC<7> B_LBLT<6> B_LBLT<7> B_LWL<6> B_XWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> A_XWL<5> B_LBLC<6> 
+ B_LBLC<5> B_LBLT<6> B_LBLT<5> B_LWL<5> B_XWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> A_XWL<4> B_LBLC<4> 
+ B_LBLC<5> B_LBLT<4> B_LBLT<5> B_LWL<4> B_XWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> A_XWL<3> B_LBLC<4> 
+ B_LBLC<3> B_LBLT<4> B_LBLT<3> B_LWL<3> B_XWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> A_XWL<2> B_LBLC<2> 
+ B_LBLC<3> B_LBLT<2> B_LBLT<3> B_LWL<2> B_XWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> A_XWL<1> B_LBLC<2> 
+ B_LBLC<1> B_LBLT<2> B_LBLT<1> B_LWL<1> B_XWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> A_XWL<0> 
+ B_BLC_BOT<0> B_LBLC<1> B_BLT_BOT<0> B_LBLT<1> B_LWL<0> B_XWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_TAP A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XIEDGEBP_COL1<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_EDGE_TB
XITAP<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_TAP
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_TAP_LR NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_TAP_LR
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX12 A Z VDD VSS
MN1 Z net6 VSS VSS sg13_lv_nmos m=1 w=4.23u l=130.00n ng=6 nrd=0 nrs=0
MN0 net6 A VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD sg13_lv_pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD sg13_lv_pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX12 A Z VDD VSS
MN1 Z net6 VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS sg13_lv_nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD sg13_lv_pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XL2<258> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<257> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<256> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<255> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<254> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<253> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<252> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<251> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<250> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<249> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<248> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<247> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<246> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<245> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<244> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<243> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<242> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<241> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<240> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<239> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<238> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<237> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<236> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<235> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<234> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<233> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<232> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<231> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<230> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<229> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<228> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<227> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<226> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<225> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<224> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<223> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<222> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<221> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<220> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<219> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<218> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<217> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<216> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<215> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<214> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<213> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<212> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<211> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<210> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<209> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<208> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<207> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<206> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<205> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<204> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<203> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<202> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<201> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<200> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<199> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<198> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<197> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<196> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<195> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<194> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<193> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<192> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<191> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<190> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<189> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<188> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<187> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<186> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<185> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<184> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<183> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<182> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<181> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<180> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<179> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<178> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<177> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<176> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<175> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<174> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<173> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_2P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net017 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net017 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net017 net8 VDD VSS / RSC_IHPSG13_CINVX2
XCAPS4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XCAPS8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI6 PULSE_L PULSE_H net017 VDD VSS / RSC_IHPSG13_XOR2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_BLDRV A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> 
+ A_SEL_P<1> A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> 
+ B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> 
+ B_SEL_P<2> B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS
MA_CWN<3> A_BLC<3> A_BLC_NMOS_DRIVE<3> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<2> A_BLC<2> A_BLC_NMOS_DRIVE<2> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<1> A_BLC<1> A_BLC_NMOS_DRIVE<1> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<0> A_BLC<0> A_BLC_NMOS_DRIVE<0> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<3> A_BLT<3> A_BLT_NMOS_DRIVE<3> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<2> A_BLT<2> A_BLT_NMOS_DRIVE<2> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<1> A_BLT<1> A_BLT_NMOS_DRIVE<1> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<0> A_BLT<0> A_BLT_NMOS_DRIVE<0> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<3> B_BLT<3> B_BLT_NMOS_DRIVE<3> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<2> B_BLT<2> B_BLT_NMOS_DRIVE<2> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<1> B_BLT<1> B_BLT_NMOS_DRIVE<1> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<0> B_BLT<0> B_BLT_NMOS_DRIVE<0> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<3> B_BLC<3> B_BLC_NMOS_DRIVE<3> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<2> B_BLC<2> B_BLC_NMOS_DRIVE<2> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<1> B_BLC<1> B_BLC_NMOS_DRIVE<1> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<0> B_BLC<0> B_BLC_NMOS_DRIVE<0> VSS VSS sg13_lv_nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CPR<3> A_BLC<3> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<2> A_BLC<2> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<1> A_BLC<1> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<0> A_BLC<0> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TWP<3> A_BLT<3> A_BLT_PMOS_DRIVE<3> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<2> A_BLT<2> A_BLT_PMOS_DRIVE<2> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<1> A_BLT<1> A_BLT_PMOS_DRIVE<1> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<0> A_BLT<0> A_BLT_PMOS_DRIVE<0> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<3> A_BLC<3> A_BLC_PMOS_DRIVE<3> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<2> A_BLC<2> A_BLC_PMOS_DRIVE<2> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<1> A_BLC<1> A_BLC_PMOS_DRIVE<1> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<0> A_BLC<0> A_BLC_PMOS_DRIVE<0> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TPR<3> A_BLT<3> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<2> A_BLT<2> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<1> A_BLT<1> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<0> A_BLT<0> A_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TSP<3> A_BLT_SEL A_SEL_N<3> A_BLT<3> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<2> A_BLT_SEL A_SEL_N<2> A_BLT<2> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<1> A_BLT_SEL A_SEL_N<1> A_BLT<1> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<0> A_BLT_SEL A_SEL_N<0> A_BLT<0> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<3> A_BLC_SEL A_SEL_N<3> A_BLC<3> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<2> A_BLC_SEL A_SEL_N<2> A_BLC<2> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<1> A_BLC_SEL A_SEL_N<1> A_BLC<1> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<0> A_BLC_SEL A_SEL_N<0> A_BLC<0> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<3> B_BLC<3> B_BLC_PMOS_DRIVE<3> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<2> B_BLC<2> B_BLC_PMOS_DRIVE<2> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<1> B_BLC<1> B_BLC_PMOS_DRIVE<1> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<0> B_BLC<0> B_BLC_PMOS_DRIVE<0> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<3> B_BLT<3> B_BLT_PMOS_DRIVE<3> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<2> B_BLT<2> B_BLT_PMOS_DRIVE<2> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<1> B_BLT<1> B_BLT_PMOS_DRIVE<1> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<0> B_BLT<0> B_BLT_PMOS_DRIVE<0> VDD VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<3> B_BLT_SEL B_SEL_N<3> B_BLT<3> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<2> B_BLT_SEL B_SEL_N<2> B_BLT<2> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<1> B_BLT_SEL B_SEL_N<1> B_BLT<1> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<0> B_BLT_SEL B_SEL_N<0> B_BLT<0> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TPR<3> B_BLT<3> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<2> B_BLT<2> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<1> B_BLT<1> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<0> B_BLT<0> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CSP<3> B_BLC_SEL B_SEL_N<3> B_BLC<3> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<2> B_BLC_SEL B_SEL_N<2> B_BLC<2> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<1> B_BLC_SEL B_SEL_N<1> B_BLC<1> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<0> B_BLC_SEL B_SEL_N<0> B_BLC<0> VDD sg13_lv_pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CPR<3> B_BLC<3> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<2> B_BLC<2> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<1> B_BLC<1> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<0> B_BLC<0> B_PRE_N VDD VDD sg13_lv_pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
XA_SEL<3> A_SEL_P<3> A_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<2> A_SEL_P<2> A_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<1> A_SEL_P<1> A_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<0> A_SEL_P<0> A_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XA_CINV<3> A_BLT_PMOS_DRIVE<3> A_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<2> A_BLT_PMOS_DRIVE<2> A_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<1> A_BLT_PMOS_DRIVE<1> A_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<0> A_BLT_PMOS_DRIVE<0> A_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<3> A_BLC_PMOS_DRIVE<3> A_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<2> A_BLC_PMOS_DRIVE<2> A_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<1> A_BLC_PMOS_DRIVE<1> A_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<0> A_BLC_PMOS_DRIVE<0> A_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_SEL<3> B_SEL_P<3> B_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<2> B_SEL_P<2> B_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<1> B_SEL_P<1> B_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<0> B_SEL_P<0> B_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XB_TINV<3> B_BLC_PMOS_DRIVE<3> B_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<2> B_BLC_PMOS_DRIVE<2> B_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<1> B_BLC_PMOS_DRIVE<1> B_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<0> B_BLC_PMOS_DRIVE<0> B_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<3> B_BLT_PMOS_DRIVE<3> B_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<2> B_BLT_PMOS_DRIVE<2> B_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<1> B_BLT_PMOS_DRIVE<1> B_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<0> B_BLT_PMOS_DRIVE<0> B_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TDEC<3> A_SEL_P<3> A_WR_ONE A_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<2> A_SEL_P<2> A_WR_ONE A_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<1> A_SEL_P<1> A_WR_ONE A_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<0> A_SEL_P<0> A_WR_ONE A_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<3> A_SEL_P<3> A_WR_ZERO A_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<2> A_SEL_P<2> A_WR_ZERO A_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<1> A_SEL_P<1> A_WR_ZERO A_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<0> A_SEL_P<0> A_WR_ZERO A_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<3> B_SEL_P<3> B_WR_ZERO B_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<2> B_SEL_P<2> B_WR_ZERO B_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<1> B_SEL_P<1> B_WR_ZERO B_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<0> B_SEL_P<0> B_WR_ZERO B_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<3> B_SEL_P<3> B_WR_ONE B_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<2> B_SEL_P<2> B_WR_ONE B_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<1> B_SEL_P<1> B_WR_ONE B_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<0> B_SEL_P<0> B_WR_ONE B_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
.ENDS
.SUBCKT RSC_IHPSG13_AND2X6 A B Z VDD VSS
MN3 Z net6 VSS VSS sg13_lv_nmos m=1 w=2.94u l=130.00n ng=3 nrd=0 nrs=0
MN4 net9 B VSS VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS sg13_lv_nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD sg13_lv_pmos m=1 w=4.86u l=130.00n ng=3 nrd=0 nrs=0
MP0 net6 B VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD sg13_lv_pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL<1> B_ADDR_COL<0> 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<31> B_BLC<30> B_BLC<29> B_BLC<28> B_BLC<27> B_BLC<26> 
+ B_BLC<25> B_BLC<24> B_BLC<23> B_BLC<22> B_BLC<21> B_BLC<20> B_BLC<19> 
+ B_BLC<18> B_BLC<17> B_BLC<16> B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> 
+ B_BLC<11> B_BLC<10> B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> 
+ B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> 
+ B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT<23> B_BLT<22> B_BLT<21> 
+ B_BLT<20> B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT<15> B_BLT<14> 
+ B_BLT<13> B_BLT<12> B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> 
+ B_BLT<5> B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L 
+ B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L 
+ B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80<1> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I80<0> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_INV<6> B_N1<1> B_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<5> B_N0<1> B_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<4> B_N0<0> B_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<3> B_ADDR_COL<1> B_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<2> B_ADDR_COL<1> B_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_ADDR_COL<0> B_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL<0> B_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<3> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<2> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<1> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL8<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XAB_BLMUX<7> A_BLC<31> A_BLC<30> A_BLC<29> A_BLC<28> A_BLC_SEL A_BLT<31> 
+ A_BLT<30> A_BLT<29> A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<31> A_SEL_P<30> 
+ A_SEL_P<29> A_SEL_P<28> A_WR_ONE A_WR_ZERO B_BLC<31> B_BLC<30> B_BLC<29> 
+ B_BLC<28> B_BLC_SEL B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> B_BLT_SEL 
+ B_PRE_N B_SEL_P<31> B_SEL_P<30> B_SEL_P<29> B_SEL_P<28> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<6> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> A_BLC_SEL A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<27> A_SEL_P<26> 
+ A_SEL_P<25> A_SEL_P<24> A_WR_ONE A_WR_ZERO B_BLC<27> B_BLC<26> B_BLC<25> 
+ B_BLC<24> B_BLC_SEL B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT_SEL 
+ B_PRE_N B_SEL_P<27> B_SEL_P<26> B_SEL_P<25> B_SEL_P<24> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<5> A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC_SEL A_BLT<23> 
+ A_BLT<22> A_BLT<21> A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<23> A_SEL_P<22> 
+ A_SEL_P<21> A_SEL_P<20> A_WR_ONE A_WR_ZERO B_BLC<23> B_BLC<22> B_BLC<21> 
+ B_BLC<20> B_BLC_SEL B_BLT<23> B_BLT<22> B_BLT<21> B_BLT<20> B_BLT_SEL 
+ B_PRE_N B_SEL_P<23> B_SEL_P<22> B_SEL_P<21> B_SEL_P<20> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<4> A_BLC<19> A_BLC<18> A_BLC<17> A_BLC<16> A_BLC_SEL A_BLT<19> 
+ A_BLT<18> A_BLT<17> A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<19> A_SEL_P<18> 
+ A_SEL_P<17> A_SEL_P<16> A_WR_ONE A_WR_ZERO B_BLC<19> B_BLC<18> B_BLC<17> 
+ B_BLC<16> B_BLC_SEL B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT_SEL 
+ B_PRE_N B_SEL_P<19> B_SEL_P<18> B_SEL_P<17> B_SEL_P<16> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_BLDRV
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<31> net041<0> B_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<30> net041<1> B_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<29> net041<2> B_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<28> net041<3> B_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<27> net041<4> B_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<26> net041<5> B_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<25> net041<6> B_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<24> net041<7> B_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<23> net041<8> B_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<22> net041<9> B_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<21> net041<10> B_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<20> net041<11> B_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<19> net041<12> B_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<18> net041<13> B_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<17> net041<14> B_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<16> net041<15> B_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net041<16> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net041<17> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net041<18> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net041<19> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net041<20> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net041<21> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net041<22> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net041<23> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net041<24> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net041<25> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net041<26> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net041<27> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net041<28> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net041<29> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net041<30> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net041<31> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net042 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DEC3<31> B_P1<1> B_P0<1> B_ADDR_DEC<7> net041<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<30> B_P1<1> B_P0<1> B_ADDR_DEC<6> net041<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<29> B_P1<1> B_P0<1> B_ADDR_DEC<5> net041<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<28> B_P1<1> B_P0<1> B_ADDR_DEC<4> net041<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<27> B_P1<1> B_P0<1> B_ADDR_DEC<3> net041<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<26> B_P1<1> B_P0<1> B_ADDR_DEC<2> net041<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<25> B_P1<1> B_P0<1> B_ADDR_DEC<1> net041<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<24> B_P1<1> B_P0<1> B_ADDR_DEC<0> net041<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<23> B_P1<1> B_N0<1> B_ADDR_DEC<7> net041<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<22> B_P1<1> B_N0<1> B_ADDR_DEC<6> net041<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<21> B_P1<1> B_N0<1> B_ADDR_DEC<5> net041<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<20> B_P1<1> B_N0<1> B_ADDR_DEC<4> net041<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<19> B_P1<1> B_N0<1> B_ADDR_DEC<3> net041<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<18> B_P1<1> B_N0<1> B_ADDR_DEC<2> net041<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<17> B_P1<1> B_N0<1> B_ADDR_DEC<1> net041<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<16> B_P1<1> B_N0<1> B_ADDR_DEC<0> net041<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<15> B_N1<0> B_P0<0> B_ADDR_DEC<7> net041<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<14> B_N1<0> B_P0<0> B_ADDR_DEC<6> net041<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<13> B_N1<0> B_P0<0> B_ADDR_DEC<5> net041<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<12> B_N1<0> B_P0<0> B_ADDR_DEC<4> net041<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<11> B_N1<0> B_P0<0> B_ADDR_DEC<3> net041<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<10> B_N1<0> B_P0<0> B_ADDR_DEC<2> net041<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<9> B_N1<0> B_P0<0> B_ADDR_DEC<1> net041<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<8> B_N1<0> B_P0<0> B_ADDR_DEC<0> net041<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<7> B_N1<0> B_N0<0> B_ADDR_DEC<7> net041<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<6> B_N1<0> B_N0<0> B_ADDR_DEC<6> net041<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<5> B_N1<0> B_N0<0> B_ADDR_DEC<5> net041<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<4> B_N1<0> B_N0<0> B_ADDR_DEC<4> net041<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<3> B_N1<0> B_N0<0> B_ADDR_DEC<3> net041<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<2> B_N1<0> B_N0<0> B_ADDR_DEC<2> net041<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<1> B_N1<0> B_N0<0> B_ADDR_DEC<1> net041<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<0> B_N1<0> B_N0<0> B_ADDR_DEC<0> net041<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4 VDD VSS
XI0<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RSC_IHPSG13_CBUFX16 A Z VDD VSS
MN0 net4 A VSS VSS sg13_lv_nmos m=1 w=2.115u l=130.00n ng=3 nrd=0 nrs=0
MN1 Z net4 VSS VSS sg13_lv_nmos m=1 w=5.64u l=130.00n ng=8 nrd=0 nrs=0
MP1 Z net4 VDD VDD sg13_lv_pmos m=1 w=13.000u l=130.00n ng=8 nrd=0 
+ nrs=0
MP0 net4 A VDD VDD sg13_lv_pmos m=1 w=4.89u l=130.00n ng=3 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX16 A Z VDD VSS
MN1 Z net6 VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS sg13_lv_nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD sg13_lv_pmos m=1 w=12.96u l=130.00n ng=8 nrd=0 nrs=0
MP0 net6 A VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1 VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI10 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> B_BLC<11> B_BLC<10> 
+ B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC<3> B_BLC<2> 
+ B_BLC<1> B_BLC<0> B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT<11> 
+ B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT<3> 
+ B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R 
+ B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L 
+ B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XI_FILL4<26> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<25> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<24> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<23> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<22> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<21> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<20> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<19> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<18> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_N0 B_P0 VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL B_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<1> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_BLDRV
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net044<0> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net044<1> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net044<2> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net044<3> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net044<4> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net044<5> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net044<6> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net044<7> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net044<8> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net044<9> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net044<10> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net044<11> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net044<12> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net044<13> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net044<14> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net044<15> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<15> B_P0 B_ADDR_DEC<7> net044<0> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<14> B_P0 B_ADDR_DEC<6> net044<1> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<13> B_P0 B_ADDR_DEC<5> net044<2> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<12> B_P0 B_ADDR_DEC<4> net044<3> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<11> B_P0 B_ADDR_DEC<3> net044<4> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<10> B_P0 B_ADDR_DEC<2> net044<5> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<9> B_P0 B_ADDR_DEC<1> net044<6> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<8> B_P0 B_ADDR_DEC<0> net044<7> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<7> B_N0 B_ADDR_DEC<7> net044<8> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<6> B_N0 B_ADDR_DEC<6> net044<9> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<5> B_N0 B_ADDR_DEC<5> net044<10> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<4> B_N0 B_ADDR_DEC<4> net044<11> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<3> B_N0 B_ADDR_DEC<3> net044<12> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<2> B_N0 B_ADDR_DEC<2> net044<13> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<1> B_N0 B_ADDR_DEC<1> net044<14> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<0> B_N0 B_ADDR_DEC<0> net044<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2P CP DN DP QN QP VDD VSS
XI_AMP CP DN DP QN QP VDD VSS / RSC_IHPSG13_DFPQD_MSAFFX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<7> B_ADDR_DEC<6> 
+ B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> 
+ B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<7> B_BLT<6> B_BLT<5> 
+ B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R 
+ B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R 
+ B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net044 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC_SEL B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I80 B_WCLK_B_L B_RCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DO_WRITE_P B_DI_N B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I75 B_DO_WRITE_P B_DI_R B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XI1<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI80<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<31> A_BLC<31> A_BLC_SEL A_BLT<31> A_BLT_SEL A_PRE_N A_SEL_P<31> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<30> A_BLC<30> A_BLC_SEL A_BLT<30> A_BLT_SEL A_PRE_N A_SEL_P<30> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<29> A_BLC<29> A_BLC_SEL A_BLT<29> A_BLT_SEL A_PRE_N A_SEL_P<29> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<28> A_BLC<28> A_BLC_SEL A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<28> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<27> A_BLC<27> A_BLC_SEL A_BLT<27> A_BLT_SEL A_PRE_N A_SEL_P<27> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<26> A_BLC<26> A_BLC_SEL A_BLT<26> A_BLT_SEL A_PRE_N A_SEL_P<26> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<25> A_BLC<25> A_BLC_SEL A_BLT<25> A_BLT_SEL A_PRE_N A_SEL_P<25> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<24> A_BLC<24> A_BLC_SEL A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<24> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<23> A_BLC<23> A_BLC_SEL A_BLT<23> A_BLT_SEL A_PRE_N A_SEL_P<23> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<22> A_BLC<22> A_BLC_SEL A_BLT<22> A_BLT_SEL A_PRE_N A_SEL_P<22> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<21> A_BLC<21> A_BLC_SEL A_BLT<21> A_BLT_SEL A_PRE_N A_SEL_P<21> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<20> A_BLC<20> A_BLC_SEL A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<20> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<19> A_BLC<19> A_BLC_SEL A_BLT<19> A_BLT_SEL A_PRE_N A_SEL_P<19> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<18> A_BLC<18> A_BLC_SEL A_BLT<18> A_BLT_SEL A_PRE_N A_SEL_P<18> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<17> A_BLC<17> A_BLC_SEL A_BLT<17> A_BLT_SEL A_PRE_N A_SEL_P<17> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<16> A_BLC<16> A_BLC_SEL A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<16> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_256x8_c2_1P_BLDRV
XA_CAPS<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS



.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX8 A Z VDD VSS
MN1 Z net6 VSS VSS sg13_lv_nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS sg13_lv_nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD sg13_lv_pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MP0 net6 A VDD VDD sg13_lv_pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> PADR<0> PADR<1> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> NADR<0> PADR<1> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> PADR<0> NADR<1> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<0> NADR<1> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI17<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI14<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI14<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI14<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI14<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<3> B_ADDR_DEC<2> 
+ B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<3> 
+ B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I 
+ B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R 
+ B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD 
+ VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I44 B_WCLK_B_L B_BM_N B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_WCLK_B_L A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XAB_BLMUX A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_256x8_c2_2P_BLDRV
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net039 net040 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I51 net039 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC03
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC01
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC02
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_2P_DEC00
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_2P_DEC04
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_2P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_TAP BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XITAP<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_1P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_256x8_c2_1P_BITKIT_TAP
XIEDGEBP_COL1<1> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_256x8_c2_1P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_256x8_c2_1P_BITKIT_TAP_LR
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0 VDD VSS / RSC_IHPSG13_FILLCAP4
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_256x8_c2_1P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC03
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC00
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC01
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_256x8_c2_1P_DEC02
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_256x8_c2_1P_DEC04
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_256x8_c2_1P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0 A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> B_BLC_BOT<1> B_BLC_BOT<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT_BOT<1> B_BLT_BOT<0> B_BLT_TOP<1> B_BLT_TOP<0> B_LWL<63> B_LWL<62> B_LWL<61> B_LWL<60> B_LWL<59> B_LWL<58> B_LWL<57> B_LWL<56> B_LWL<55> B_LWL<54> B_LWL<53> B_LWL<52> B_LWL<51> B_LWL<50> B_LWL<49> B_LWL<48> B_LWL<47> B_LWL<46> B_LWL<45> B_LWL<44> B_LWL<43> B_LWL<42> B_LWL<41> B_LWL<40> B_LWL<39> B_LWL<38> B_LWL<37> B_LWL<36> B_LWL<35> B_LWL<34> B_LWL<33> B_LWL<32> B_LWL<31> B_LWL<30> B_LWL<29> B_LWL<28> B_LWL<27> B_LWL<26> B_LWL<25> B_LWL<24> B_LWL<23> B_LWL<22> B_LWL<21> B_LWL<20> B_LWL<19> B_LWL<18> B_LWL<17> B_LWL<16> B_LWL<15> B_LWL<14> B_LWL<13> B_LWL<12> B_LWL<11> B_LWL<10> B_LWL<9> B_LWL<8> B_LWL<7> B_LWL<6> B_LWL<5> B_LWL<4> B_LWL<3> B_LWL<2> B_LWL<1> B_LWL<0> B_RWL<63> B_RWL<62> B_RWL<61> B_RWL<60> B_RWL<59> B_RWL<58> B_RWL<57> B_RWL<56> B_RWL<55> B_RWL<54> B_RWL<53> B_RWL<52> B_RWL<51> B_RWL<50> B_RWL<49> B_RWL<48> B_RWL<47> B_RWL<46> B_RWL<45> B_RWL<44> B_RWL<43> B_RWL<42> B_RWL<41> B_RWL<40> B_RWL<39> B_RWL<38> B_RWL<37> B_RWL<36> B_RWL<35> B_RWL<34> B_RWL<33> B_RWL<32> B_RWL<31> B_RWL<30> B_RWL<29> B_RWL<28> B_RWL<27> B_RWL<26> B_RWL<25> B_RWL<24> B_RWL<23> B_RWL<22> B_RWL<21> B_RWL<20> B_RWL<19> B_RWL<18> B_RWL<17> B_RWL<16> B_RWL<15> B_RWL<14> B_RWL<13> B_RWL<12> B_RWL<11> B_RWL<10> B_RWL<9> B_RWL<8> B_RWL<7> B_RWL<6> B_RWL<5> B_RWL<4> B_RWL<3> B_RWL<2> B_RWL<1> B_RWL<0> VDD_CORE VSS
XRAM<4> A_BLC<5> A_BLC<4> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<5> A_BLT<4> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> B_BLC<5> B_BLC<4> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT<5> B_BLT<4> B_BLT_TOP<1> B_BLT_TOP<0> B_LWL<63> B_LWL<62> B_LWL<61> B_LWL<60> B_LWL<59> B_LWL<58> B_LWL<57> B_LWL<56> B_LWL<55> B_LWL<54> B_LWL<53> B_LWL<52> B_LWL<51> B_LWL<50> B_LWL<49> B_LWL<48> B_RWL<63> B_RWL<62> B_RWL<61> B_RWL<60> B_RWL<59> B_RWL<58> B_RWL<57> B_RWL<56> B_RWL<55> B_RWL<54> B_RWL<53> B_RWL<52> B_RWL<51> B_RWL<50> B_RWL<49> B_RWL<48> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_SRAM
XRAM<3> A_BLC<3> A_BLC<2> A_BLC<5> A_BLC<4> A_BLT<3> A_BLT<2> A_BLT<5> A_BLT<4> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> B_BLC<3> B_BLC<2> B_BLC<5> B_BLC<4> B_BLT<3> B_BLT<2> B_BLT<5> B_BLT<4> B_LWL<47> B_LWL<46> B_LWL<45> B_LWL<44> B_LWL<43> B_LWL<42> B_LWL<41> B_LWL<40> B_LWL<39> B_LWL<38> B_LWL<37> B_LWL<36> B_LWL<35> B_LWL<34> B_LWL<33> B_LWL<32> B_RWL<47> B_RWL<46> B_RWL<45> B_RWL<44> B_RWL<43> B_RWL<42> B_RWL<41> B_RWL<40> B_RWL<39> B_RWL<38> B_RWL<37> B_RWL<36> B_RWL<35> B_RWL<34> B_RWL<33> B_RWL<32> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_SRAM
XRAM<2> A_BLC<1> A_BLC<0> A_BLC<3> A_BLC<2> A_BLT<1> A_BLT<0> A_BLT<3> A_BLT<2> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> B_BLC<1> B_BLC<0> B_BLC<3> B_BLC<2> B_BLT<1> B_BLT<0> B_BLT<3> B_BLT<2> B_LWL<31> B_LWL<30> B_LWL<29> B_LWL<28> B_LWL<27> B_LWL<26> B_LWL<25> B_LWL<24> B_LWL<23> B_LWL<22> B_LWL<21> B_LWL<20> B_LWL<19> B_LWL<18> B_LWL<17> B_LWL<16> B_RWL<31> B_RWL<30> B_RWL<29> B_RWL<28> B_RWL<27> B_RWL<26> B_RWL<25> B_RWL<24> B_RWL<23> B_RWL<22> B_RWL<21> B_RWL<20> B_RWL<19> B_RWL<18> B_RWL<17> B_RWL<16> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_SRAM
XRAM<1> A_BLC_BOT<1> A_BLC_BOT<0> A_BLC<1> A_BLC<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT<1> A_BLT<0> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> B_BLC_BOT<1> B_BLC_BOT<0> B_BLC<1> B_BLC<0> B_BLT_BOT<1> B_BLT_BOT<0> B_BLT<1> B_BLT<0> B_LWL<15> B_LWL<14> B_LWL<13> B_LWL<12> B_LWL<11> B_LWL<10> B_LWL<9> B_LWL<8> B_LWL<7> B_LWL<6> B_LWL<5> B_LWL<4> B_LWL<3> B_LWL<2> B_LWL<1> B_LWL<0> B_RWL<15> B_RWL<14> B_RWL<13> B_RWL<12> B_RWL<11> B_RWL<10> B_RWL<9> B_RWL<8> B_RWL<7> B_RWL<6> B_RWL<5> B_RWL<4> B_RWL<3> B_RWL<2> B_RWL<1> B_RWL<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_SRAM
XEDGE<1> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_TOP<1> A_BLT_TOP<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT_TOP<1> B_BLT_TOP<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_TB
XEDGE<0> A_BLC_BOT<1> A_BLC_BOT<0> A_BLT_BOT<1> A_BLT_BOT<0> B_BLC_BOT<1> B_BLC_BOT<0> B_BLT_BOT<1> B_BLT_BOT<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_TB
.ENDS




.SUBCKT RM_IHPSG13_256x8_c2_2P_MATRIX_pcell_1 A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> B_BLC<11> B_BLC<10> B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_WL<63> B_WL<62> B_WL<61> B_WL<60> B_WL<59> B_WL<58> B_WL<57> B_WL<56> B_WL<55> B_WL<54> B_WL<53> B_WL<52> B_WL<51> B_WL<50> B_WL<49> B_WL<48> B_WL<47> B_WL<46> B_WL<45> B_WL<44> B_WL<43> B_WL<42> B_WL<41> B_WL<40> B_WL<39> B_WL<38> B_WL<37> B_WL<36> B_WL<35> B_WL<34> B_WL<33> B_WL<32> B_WL<31> B_WL<30> B_WL<29> B_WL<28> B_WL<27> B_WL<26> B_WL<25> B_WL<24> B_WL<23> B_WL<22> B_WL<21> B_WL<20> B_WL<19> B_WL<18> B_WL<17> B_WL<16> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> B_WL<1> B_WL<0> VDD_CORE VSS
XCORNER<3> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_CORNER
XCORNER<2> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_CORNER
XCORNER<1> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_CORNER
XCORNER<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_CORNER
XRAMEDGE_L<3> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> B_WL<63> B_WL<62> B_WL<61> B_WL<60> B_WL<59> B_WL<58> B_WL<57> B_WL<56> B_WL<55> B_WL<54> B_WL<53> B_WL<52> B_WL<51> B_WL<50> B_WL<49> B_WL<48> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<2> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> B_WL<47> B_WL<46> B_WL<45> B_WL<44> B_WL<43> B_WL<42> B_WL<41> B_WL<40> B_WL<39> B_WL<38> B_WL<37> B_WL<36> B_WL<35> B_WL<34> B_WL<33> B_WL<32> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<1> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> B_WL<31> B_WL<30> B_WL<29> B_WL<28> B_WL<27> B_WL<26> B_WL<25> B_WL<24> B_WL<23> B_WL<22> B_WL<21> B_WL<20> B_WL<19> B_WL<18> B_WL<17> B_WL<16> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<0> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> B_WL<1> B_WL<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<3> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> B_IWL<511> B_IWL<510> B_IWL<509> B_IWL<508> B_IWL<507> B_IWL<506> B_IWL<505> B_IWL<504> B_IWL<503> B_IWL<502> B_IWL<501> B_IWL<500> B_IWL<499> B_IWL<498> B_IWL<497> B_IWL<496> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<2> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> B_IWL<495> B_IWL<494> B_IWL<493> B_IWL<492> B_IWL<491> B_IWL<490> B_IWL<489> B_IWL<488> B_IWL<487> B_IWL<486> B_IWL<485> B_IWL<484> B_IWL<483> B_IWL<482> B_IWL<481> B_IWL<480> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<1> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> B_IWL<479> B_IWL<478> B_IWL<477> B_IWL<476> B_IWL<475> B_IWL<474> B_IWL<473> B_IWL<472> B_IWL<471> B_IWL<470> B_IWL<469> B_IWL<468> B_IWL<467> B_IWL<466> B_IWL<465> B_IWL<464> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<0> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> B_IWL<463> B_IWL<462> B_IWL<461> B_IWL<460> B_IWL<459> B_IWL<458> B_IWL<457> B_IWL<456> B_IWL<455> B_IWL<454> B_IWL<453> B_IWL<452> B_IWL<451> B_IWL<450> B_IWL<449> B_IWL<448> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_BITKIT_16x2_EDGE_LR
XCOL<7> A_BLC<15> A_BLC<14> A_BLC_TOP<15> A_BLC_TOP<14> A_BLT<15> A_BLT<14> A_BLT_TOP<15> A_BLT_TOP<14> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> B_BLC<15> B_BLC<14> B_BLC_TOP<15> B_BLC_TOP<14> B_BLT<15> B_BLT<14> B_BLT_TOP<15> B_BLT_TOP<14> B_IWL<447> B_IWL<446> B_IWL<445> B_IWL<444> B_IWL<443> B_IWL<442> B_IWL<441> B_IWL<440> B_IWL<439> B_IWL<438> B_IWL<437> B_IWL<436> B_IWL<435> B_IWL<434> B_IWL<433> B_IWL<432> B_IWL<431> B_IWL<430> B_IWL<429> B_IWL<428> B_IWL<427> B_IWL<426> B_IWL<425> B_IWL<424> B_IWL<423> B_IWL<422> B_IWL<421> B_IWL<420> B_IWL<419> B_IWL<418> B_IWL<417> B_IWL<416> B_IWL<415> B_IWL<414> B_IWL<413> B_IWL<412> B_IWL<411> B_IWL<410> B_IWL<409> B_IWL<408> B_IWL<407> B_IWL<406> B_IWL<405> B_IWL<404> B_IWL<403> B_IWL<402> B_IWL<401> B_IWL<400> B_IWL<399> B_IWL<398> B_IWL<397> B_IWL<396> B_IWL<395> B_IWL<394> B_IWL<393> B_IWL<392> B_IWL<391> B_IWL<390> B_IWL<389> B_IWL<388> B_IWL<387> B_IWL<386> B_IWL<385> B_IWL<384> B_IWL<511> B_IWL<510> B_IWL<509> B_IWL<508> B_IWL<507> B_IWL<506> B_IWL<505> B_IWL<504> B_IWL<503> B_IWL<502> B_IWL<501> B_IWL<500> B_IWL<499> B_IWL<498> B_IWL<497> B_IWL<496> B_IWL<495> B_IWL<494> B_IWL<493> B_IWL<492> B_IWL<491> B_IWL<490> B_IWL<489> B_IWL<488> B_IWL<487> B_IWL<486> B_IWL<485> B_IWL<484> B_IWL<483> B_IWL<482> B_IWL<481> B_IWL<480> B_IWL<479> B_IWL<478> B_IWL<477> B_IWL<476> B_IWL<475> B_IWL<474> B_IWL<473> B_IWL<472> B_IWL<471> B_IWL<470> B_IWL<469> B_IWL<468> B_IWL<467> B_IWL<466> B_IWL<465> B_IWL<464> B_IWL<463> B_IWL<462> B_IWL<461> B_IWL<460> B_IWL<459> B_IWL<458> B_IWL<457> B_IWL<456> B_IWL<455> B_IWL<454> B_IWL<453> B_IWL<452> B_IWL<451> B_IWL<450> B_IWL<449> B_IWL<448> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<6> A_BLC<13> A_BLC<12> A_BLC_TOP<13> A_BLC_TOP<12> A_BLT<13> A_BLT<12> A_BLT_TOP<13> A_BLT_TOP<12> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> B_BLC<13> B_BLC<12> B_BLC_TOP<13> B_BLC_TOP<12> B_BLT<13> B_BLT<12> B_BLT_TOP<13> B_BLT_TOP<12> B_IWL<383> B_IWL<382> B_IWL<381> B_IWL<380> B_IWL<379> B_IWL<378> B_IWL<377> B_IWL<376> B_IWL<375> B_IWL<374> B_IWL<373> B_IWL<372> B_IWL<371> B_IWL<370> B_IWL<369> B_IWL<368> B_IWL<367> B_IWL<366> B_IWL<365> B_IWL<364> B_IWL<363> B_IWL<362> B_IWL<361> B_IWL<360> B_IWL<359> B_IWL<358> B_IWL<357> B_IWL<356> B_IWL<355> B_IWL<354> B_IWL<353> B_IWL<352> B_IWL<351> B_IWL<350> B_IWL<349> B_IWL<348> B_IWL<347> B_IWL<346> B_IWL<345> B_IWL<344> B_IWL<343> B_IWL<342> B_IWL<341> B_IWL<340> B_IWL<339> B_IWL<338> B_IWL<337> B_IWL<336> B_IWL<335> B_IWL<334> B_IWL<333> B_IWL<332> B_IWL<331> B_IWL<330> B_IWL<329> B_IWL<328> B_IWL<327> B_IWL<326> B_IWL<325> B_IWL<324> B_IWL<323> B_IWL<322> B_IWL<321> B_IWL<320> B_IWL<447> B_IWL<446> B_IWL<445> B_IWL<444> B_IWL<443> B_IWL<442> B_IWL<441> B_IWL<440> B_IWL<439> B_IWL<438> B_IWL<437> B_IWL<436> B_IWL<435> B_IWL<434> B_IWL<433> B_IWL<432> B_IWL<431> B_IWL<430> B_IWL<429> B_IWL<428> B_IWL<427> B_IWL<426> B_IWL<425> B_IWL<424> B_IWL<423> B_IWL<422> B_IWL<421> B_IWL<420> B_IWL<419> B_IWL<418> B_IWL<417> B_IWL<416> B_IWL<415> B_IWL<414> B_IWL<413> B_IWL<412> B_IWL<411> B_IWL<410> B_IWL<409> B_IWL<408> B_IWL<407> B_IWL<406> B_IWL<405> B_IWL<404> B_IWL<403> B_IWL<402> B_IWL<401> B_IWL<400> B_IWL<399> B_IWL<398> B_IWL<397> B_IWL<396> B_IWL<395> B_IWL<394> B_IWL<393> B_IWL<392> B_IWL<391> B_IWL<390> B_IWL<389> B_IWL<388> B_IWL<387> B_IWL<386> B_IWL<385> B_IWL<384> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<5> A_BLC<11> A_BLC<10> A_BLC_TOP<11> A_BLC_TOP<10> A_BLT<11> A_BLT<10> A_BLT_TOP<11> A_BLT_TOP<10> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> B_BLC<11> B_BLC<10> B_BLC_TOP<11> B_BLC_TOP<10> B_BLT<11> B_BLT<10> B_BLT_TOP<11> B_BLT_TOP<10> B_IWL<319> B_IWL<318> B_IWL<317> B_IWL<316> B_IWL<315> B_IWL<314> B_IWL<313> B_IWL<312> B_IWL<311> B_IWL<310> B_IWL<309> B_IWL<308> B_IWL<307> B_IWL<306> B_IWL<305> B_IWL<304> B_IWL<303> B_IWL<302> B_IWL<301> B_IWL<300> B_IWL<299> B_IWL<298> B_IWL<297> B_IWL<296> B_IWL<295> B_IWL<294> B_IWL<293> B_IWL<292> B_IWL<291> B_IWL<290> B_IWL<289> B_IWL<288> B_IWL<287> B_IWL<286> B_IWL<285> B_IWL<284> B_IWL<283> B_IWL<282> B_IWL<281> B_IWL<280> B_IWL<279> B_IWL<278> B_IWL<277> B_IWL<276> B_IWL<275> B_IWL<274> B_IWL<273> B_IWL<272> B_IWL<271> B_IWL<270> B_IWL<269> B_IWL<268> B_IWL<267> B_IWL<266> B_IWL<265> B_IWL<264> B_IWL<263> B_IWL<262> B_IWL<261> B_IWL<260> B_IWL<259> B_IWL<258> B_IWL<257> B_IWL<256> B_IWL<383> B_IWL<382> B_IWL<381> B_IWL<380> B_IWL<379> B_IWL<378> B_IWL<377> B_IWL<376> B_IWL<375> B_IWL<374> B_IWL<373> B_IWL<372> B_IWL<371> B_IWL<370> B_IWL<369> B_IWL<368> B_IWL<367> B_IWL<366> B_IWL<365> B_IWL<364> B_IWL<363> B_IWL<362> B_IWL<361> B_IWL<360> B_IWL<359> B_IWL<358> B_IWL<357> B_IWL<356> B_IWL<355> B_IWL<354> B_IWL<353> B_IWL<352> B_IWL<351> B_IWL<350> B_IWL<349> B_IWL<348> B_IWL<347> B_IWL<346> B_IWL<345> B_IWL<344> B_IWL<343> B_IWL<342> B_IWL<341> B_IWL<340> B_IWL<339> B_IWL<338> B_IWL<337> B_IWL<336> B_IWL<335> B_IWL<334> B_IWL<333> B_IWL<332> B_IWL<331> B_IWL<330> B_IWL<329> B_IWL<328> B_IWL<327> B_IWL<326> B_IWL<325> B_IWL<324> B_IWL<323> B_IWL<322> B_IWL<321> B_IWL<320> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<4> A_BLC<9> A_BLC<8> A_BLC_TOP<9> A_BLC_TOP<8> A_BLT<9> A_BLT<8> A_BLT_TOP<9> A_BLT_TOP<8> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> B_BLC<9> B_BLC<8> B_BLC_TOP<9> B_BLC_TOP<8> B_BLT<9> B_BLT<8> B_BLT_TOP<9> B_BLT_TOP<8> B_IWL<255> B_IWL<254> B_IWL<253> B_IWL<252> B_IWL<251> B_IWL<250> B_IWL<249> B_IWL<248> B_IWL<247> B_IWL<246> B_IWL<245> B_IWL<244> B_IWL<243> B_IWL<242> B_IWL<241> B_IWL<240> B_IWL<239> B_IWL<238> B_IWL<237> B_IWL<236> B_IWL<235> B_IWL<234> B_IWL<233> B_IWL<232> B_IWL<231> B_IWL<230> B_IWL<229> B_IWL<228> B_IWL<227> B_IWL<226> B_IWL<225> B_IWL<224> B_IWL<223> B_IWL<222> B_IWL<221> B_IWL<220> B_IWL<219> B_IWL<218> B_IWL<217> B_IWL<216> B_IWL<215> B_IWL<214> B_IWL<213> B_IWL<212> B_IWL<211> B_IWL<210> B_IWL<209> B_IWL<208> B_IWL<207> B_IWL<206> B_IWL<205> B_IWL<204> B_IWL<203> B_IWL<202> B_IWL<201> B_IWL<200> B_IWL<199> B_IWL<198> B_IWL<197> B_IWL<196> B_IWL<195> B_IWL<194> B_IWL<193> B_IWL<192> B_IWL<319> B_IWL<318> B_IWL<317> B_IWL<316> B_IWL<315> B_IWL<314> B_IWL<313> B_IWL<312> B_IWL<311> B_IWL<310> B_IWL<309> B_IWL<308> B_IWL<307> B_IWL<306> B_IWL<305> B_IWL<304> B_IWL<303> B_IWL<302> B_IWL<301> B_IWL<300> B_IWL<299> B_IWL<298> B_IWL<297> B_IWL<296> B_IWL<295> B_IWL<294> B_IWL<293> B_IWL<292> B_IWL<291> B_IWL<290> B_IWL<289> B_IWL<288> B_IWL<287> B_IWL<286> B_IWL<285> B_IWL<284> B_IWL<283> B_IWL<282> B_IWL<281> B_IWL<280> B_IWL<279> B_IWL<278> B_IWL<277> B_IWL<276> B_IWL<275> B_IWL<274> B_IWL<273> B_IWL<272> B_IWL<271> B_IWL<270> B_IWL<269> B_IWL<268> B_IWL<267> B_IWL<266> B_IWL<265> B_IWL<264> B_IWL<263> B_IWL<262> B_IWL<261> B_IWL<260> B_IWL<259> B_IWL<258> B_IWL<257> B_IWL<256> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<3> A_BLC<7> A_BLC<6> A_BLC_TOP<7> A_BLC_TOP<6> A_BLT<7> A_BLT<6> A_BLT_TOP<7> A_BLT_TOP<6> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> B_BLC<7> B_BLC<6> B_BLC_TOP<7> B_BLC_TOP<6> B_BLT<7> B_BLT<6> B_BLT_TOP<7> B_BLT_TOP<6> B_IWL<191> B_IWL<190> B_IWL<189> B_IWL<188> B_IWL<187> B_IWL<186> B_IWL<185> B_IWL<184> B_IWL<183> B_IWL<182> B_IWL<181> B_IWL<180> B_IWL<179> B_IWL<178> B_IWL<177> B_IWL<176> B_IWL<175> B_IWL<174> B_IWL<173> B_IWL<172> B_IWL<171> B_IWL<170> B_IWL<169> B_IWL<168> B_IWL<167> B_IWL<166> B_IWL<165> B_IWL<164> B_IWL<163> B_IWL<162> B_IWL<161> B_IWL<160> B_IWL<159> B_IWL<158> B_IWL<157> B_IWL<156> B_IWL<155> B_IWL<154> B_IWL<153> B_IWL<152> B_IWL<151> B_IWL<150> B_IWL<149> B_IWL<148> B_IWL<147> B_IWL<146> B_IWL<145> B_IWL<144> B_IWL<143> B_IWL<142> B_IWL<141> B_IWL<140> B_IWL<139> B_IWL<138> B_IWL<137> B_IWL<136> B_IWL<135> B_IWL<134> B_IWL<133> B_IWL<132> B_IWL<131> B_IWL<130> B_IWL<129> B_IWL<128> B_IWL<255> B_IWL<254> B_IWL<253> B_IWL<252> B_IWL<251> B_IWL<250> B_IWL<249> B_IWL<248> B_IWL<247> B_IWL<246> B_IWL<245> B_IWL<244> B_IWL<243> B_IWL<242> B_IWL<241> B_IWL<240> B_IWL<239> B_IWL<238> B_IWL<237> B_IWL<236> B_IWL<235> B_IWL<234> B_IWL<233> B_IWL<232> B_IWL<231> B_IWL<230> B_IWL<229> B_IWL<228> B_IWL<227> B_IWL<226> B_IWL<225> B_IWL<224> B_IWL<223> B_IWL<222> B_IWL<221> B_IWL<220> B_IWL<219> B_IWL<218> B_IWL<217> B_IWL<216> B_IWL<215> B_IWL<214> B_IWL<213> B_IWL<212> B_IWL<211> B_IWL<210> B_IWL<209> B_IWL<208> B_IWL<207> B_IWL<206> B_IWL<205> B_IWL<204> B_IWL<203> B_IWL<202> B_IWL<201> B_IWL<200> B_IWL<199> B_IWL<198> B_IWL<197> B_IWL<196> B_IWL<195> B_IWL<194> B_IWL<193> B_IWL<192> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<2> A_BLC<5> A_BLC<4> A_BLC_TOP<5> A_BLC_TOP<4> A_BLT<5> A_BLT<4> A_BLT_TOP<5> A_BLT_TOP<4> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> B_BLC<5> B_BLC<4> B_BLC_TOP<5> B_BLC_TOP<4> B_BLT<5> B_BLT<4> B_BLT_TOP<5> B_BLT_TOP<4> B_IWL<127> B_IWL<126> B_IWL<125> B_IWL<124> B_IWL<123> B_IWL<122> B_IWL<121> B_IWL<120> B_IWL<119> B_IWL<118> B_IWL<117> B_IWL<116> B_IWL<115> B_IWL<114> B_IWL<113> B_IWL<112> B_IWL<111> B_IWL<110> B_IWL<109> B_IWL<108> B_IWL<107> B_IWL<106> B_IWL<105> B_IWL<104> B_IWL<103> B_IWL<102> B_IWL<101> B_IWL<100> B_IWL<99> B_IWL<98> B_IWL<97> B_IWL<96> B_IWL<95> B_IWL<94> B_IWL<93> B_IWL<92> B_IWL<91> B_IWL<90> B_IWL<89> B_IWL<88> B_IWL<87> B_IWL<86> B_IWL<85> B_IWL<84> B_IWL<83> B_IWL<82> B_IWL<81> B_IWL<80> B_IWL<79> B_IWL<78> B_IWL<77> B_IWL<76> B_IWL<75> B_IWL<74> B_IWL<73> B_IWL<72> B_IWL<71> B_IWL<70> B_IWL<69> B_IWL<68> B_IWL<67> B_IWL<66> B_IWL<65> B_IWL<64> B_IWL<191> B_IWL<190> B_IWL<189> B_IWL<188> B_IWL<187> B_IWL<186> B_IWL<185> B_IWL<184> B_IWL<183> B_IWL<182> B_IWL<181> B_IWL<180> B_IWL<179> B_IWL<178> B_IWL<177> B_IWL<176> B_IWL<175> B_IWL<174> B_IWL<173> B_IWL<172> B_IWL<171> B_IWL<170> B_IWL<169> B_IWL<168> B_IWL<167> B_IWL<166> B_IWL<165> B_IWL<164> B_IWL<163> B_IWL<162> B_IWL<161> B_IWL<160> B_IWL<159> B_IWL<158> B_IWL<157> B_IWL<156> B_IWL<155> B_IWL<154> B_IWL<153> B_IWL<152> B_IWL<151> B_IWL<150> B_IWL<149> B_IWL<148> B_IWL<147> B_IWL<146> B_IWL<145> B_IWL<144> B_IWL<143> B_IWL<142> B_IWL<141> B_IWL<140> B_IWL<139> B_IWL<138> B_IWL<137> B_IWL<136> B_IWL<135> B_IWL<134> B_IWL<133> B_IWL<132> B_IWL<131> B_IWL<130> B_IWL<129> B_IWL<128> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<1> A_BLC<3> A_BLC<2> A_BLC_TOP<3> A_BLC_TOP<2> A_BLT<3> A_BLT<2> A_BLT_TOP<3> A_BLT_TOP<2> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> B_BLC<3> B_BLC<2> B_BLC_TOP<3> B_BLC_TOP<2> B_BLT<3> B_BLT<2> B_BLT_TOP<3> B_BLT_TOP<2> B_IWL<63> B_IWL<62> B_IWL<61> B_IWL<60> B_IWL<59> B_IWL<58> B_IWL<57> B_IWL<56> B_IWL<55> B_IWL<54> B_IWL<53> B_IWL<52> B_IWL<51> B_IWL<50> B_IWL<49> B_IWL<48> B_IWL<47> B_IWL<46> B_IWL<45> B_IWL<44> B_IWL<43> B_IWL<42> B_IWL<41> B_IWL<40> B_IWL<39> B_IWL<38> B_IWL<37> B_IWL<36> B_IWL<35> B_IWL<34> B_IWL<33> B_IWL<32> B_IWL<31> B_IWL<30> B_IWL<29> B_IWL<28> B_IWL<27> B_IWL<26> B_IWL<25> B_IWL<24> B_IWL<23> B_IWL<22> B_IWL<21> B_IWL<20> B_IWL<19> B_IWL<18> B_IWL<17> B_IWL<16> B_IWL<15> B_IWL<14> B_IWL<13> B_IWL<12> B_IWL<11> B_IWL<10> B_IWL<9> B_IWL<8> B_IWL<7> B_IWL<6> B_IWL<5> B_IWL<4> B_IWL<3> B_IWL<2> B_IWL<1> B_IWL<0> B_IWL<127> B_IWL<126> B_IWL<125> B_IWL<124> B_IWL<123> B_IWL<122> B_IWL<121> B_IWL<120> B_IWL<119> B_IWL<118> B_IWL<117> B_IWL<116> B_IWL<115> B_IWL<114> B_IWL<113> B_IWL<112> B_IWL<111> B_IWL<110> B_IWL<109> B_IWL<108> B_IWL<107> B_IWL<106> B_IWL<105> B_IWL<104> B_IWL<103> B_IWL<102> B_IWL<101> B_IWL<100> B_IWL<99> B_IWL<98> B_IWL<97> B_IWL<96> B_IWL<95> B_IWL<94> B_IWL<93> B_IWL<92> B_IWL<91> B_IWL<90> B_IWL<89> B_IWL<88> B_IWL<87> B_IWL<86> B_IWL<85> B_IWL<84> B_IWL<83> B_IWL<82> B_IWL<81> B_IWL<80> B_IWL<79> B_IWL<78> B_IWL<77> B_IWL<76> B_IWL<75> B_IWL<74> B_IWL<73> B_IWL<72> B_IWL<71> B_IWL<70> B_IWL<69> B_IWL<68> B_IWL<67> B_IWL<66> B_IWL<65> B_IWL<64> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
XCOL<0> A_BLC<1> A_BLC<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<1> A_BLT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> B_BLC<1> B_BLC<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT<1> B_BLT<0> B_BLT_TOP<1> B_BLT_TOP<0> B_WL<63> B_WL<62> B_WL<61> B_WL<60> B_WL<59> B_WL<58> B_WL<57> B_WL<56> B_WL<55> B_WL<54> B_WL<53> B_WL<52> B_WL<51> B_WL<50> B_WL<49> B_WL<48> B_WL<47> B_WL<46> B_WL<45> B_WL<44> B_WL<43> B_WL<42> B_WL<41> B_WL<40> B_WL<39> B_WL<38> B_WL<37> B_WL<36> B_WL<35> B_WL<34> B_WL<33> B_WL<32> B_WL<31> B_WL<30> B_WL<29> B_WL<28> B_WL<27> B_WL<26> B_WL<25> B_WL<24> B_WL<23> B_WL<22> B_WL<21> B_WL<20> B_WL<19> B_WL<18> B_WL<17> B_WL<16> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> B_WL<1> B_WL<0> B_IWL<63> B_IWL<62> B_IWL<61> B_IWL<60> B_IWL<59> B_IWL<58> B_IWL<57> B_IWL<56> B_IWL<55> B_IWL<54> B_IWL<53> B_IWL<52> B_IWL<51> B_IWL<50> B_IWL<49> B_IWL<48> B_IWL<47> B_IWL<46> B_IWL<45> B_IWL<44> B_IWL<43> B_IWL<42> B_IWL<41> B_IWL<40> B_IWL<39> B_IWL<38> B_IWL<37> B_IWL<36> B_IWL<35> B_IWL<34> B_IWL<33> B_IWL<32> B_IWL<31> B_IWL<30> B_IWL<29> B_IWL<28> B_IWL<27> B_IWL<26> B_IWL<25> B_IWL<24> B_IWL<23> B_IWL<22> B_IWL<21> B_IWL<20> B_IWL<19> B_IWL<18> B_IWL<17> B_IWL<16> B_IWL<15> B_IWL<14> B_IWL<13> B_IWL<12> B_IWL<11> B_IWL<10> B_IWL<9> B_IWL<8> B_IWL<7> B_IWL<6> B_IWL<5> B_IWL<4> B_IWL<3> B_IWL<2> B_IWL<1> B_IWL<0> VDD_CORE VSS / RM_IHPSG13_256x8_c2_2P_COLUMN_pcell_0
.ENDS




.SUBCKT RM_IHPSG13_256x8_c2_2P_DLY_pcell_2 A Z VDD VSS
	XIDL D<9> Z VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDM<9> D<8> D<9> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<8> D<7> D<8> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<7> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<6> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<5> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<4> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS


.SUBCKT RM_IHPSG13_256x8_c2_2P_DLY_pcell_3 A Z VDD VSS
	XIDM<10> D<9> Z VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<9> D<8> D<9> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<8> D<7> D<8> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<7> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<6> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<5> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<4> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS



.SUBCKT RM_IHPSG13_2P_256x8_c2_bm_bist A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> A_ADDR<1> A_ADDR<0> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_BM<7> A_BIST_BM<6> A_BIST_BM<5> A_BIST_BM<4> A_BIST_BM<3> A_BIST_BM<2> A_BIST_BM<1> A_BIST_BM<0> A_BIST_CLK A_BIST_DIN<7> A_BIST_DIN<6> A_BIST_DIN<5> A_BIST_DIN<4> A_BIST_DIN<3> A_BIST_DIN<2> A_BIST_DIN<1> A_BIST_DIN<0> A_BIST_EN A_BIST_MEN A_BIST_REN A_BIST_WEN A_BM<7> A_BM<6> A_BM<5> A_BM<4> A_BM<3> A_BM<2> A_BM<1> A_BM<0> A_CLK A_DIN<7> A_DIN<6> A_DIN<5> A_DIN<4> A_DIN<3> A_DIN<2> A_DIN<1> A_DIN<0> A_DLY A_DOUT<7> A_DOUT<6> A_DOUT<5> A_DOUT<4> A_DOUT<3> A_DOUT<2> A_DOUT<1> A_DOUT<0> A_MEN A_REN A_WEN B_ADDR<7> B_ADDR<6> B_ADDR<5> B_ADDR<4> B_ADDR<3> B_ADDR<2> B_ADDR<1> B_ADDR<0> B_BIST_ADDR<7> B_BIST_ADDR<6> B_BIST_ADDR<5> B_BIST_ADDR<4> B_BIST_ADDR<3> B_BIST_ADDR<2> B_BIST_ADDR<1> B_BIST_ADDR<0> B_BIST_BM<7> B_BIST_BM<6> B_BIST_BM<5> B_BIST_BM<4> B_BIST_BM<3> B_BIST_BM<2> B_BIST_BM<1> B_BIST_BM<0> B_BIST_CLK B_BIST_DIN<7> B_BIST_DIN<6> B_BIST_DIN<5> B_BIST_DIN<4> B_BIST_DIN<3> B_BIST_DIN<2> B_BIST_DIN<1> B_BIST_DIN<0> B_BIST_EN B_BIST_MEN B_BIST_REN B_BIST_WEN B_BM<7> B_BM<6> B_BM<5> B_BM<4> B_BM<3> B_BM<2> B_BM<1> B_BM<0> B_CLK B_DIN<7> B_DIN<6> B_DIN<5> B_DIN<4> B_DIN<3> B_DIN<2> B_DIN<1> B_DIN<0> B_DLY B_DOUT<7> B_DOUT<6> B_DOUT<5> B_DOUT<4> B_DOUT<3> B_DOUT<2> B_DOUT<1> B_DOUT<0> B_MEN B_REN B_WEN VDD! VDDARRAY! VSS!


XRAM<1> a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0> b_blc_r<15> b_blc_r<14> b_blc_r<13> b_blc_r<12> b_blc_r<11> b_blc_r<10> b_blc_r<9> b_blc_r<8> b_blc_r<7> b_blc_r<6> b_blc_r<5> b_blc_r<4> b_blc_r<3> b_blc_r<2> b_blc_r<1> b_blc_r<0> b_blt_r<15> b_blt_r<14> b_blt_r<13> b_blt_r<12> b_blt_r<11> b_blt_r<10> b_blt_r<9> b_blt_r<8> b_blt_r<7> b_blt_r<6> b_blt_r<5> b_blt_r<4> b_blt_r<3> b_blt_r<2> b_blt_r<1> b_blt_r<0> b_wl_r<63> b_wl_r<62> b_wl_r<61> b_wl_r<60> b_wl_r<59> b_wl_r<58> b_wl_r<57> b_wl_r<56> b_wl_r<55> b_wl_r<54> b_wl_r<53> b_wl_r<52> b_wl_r<51> b_wl_r<50> b_wl_r<49> b_wl_r<48> b_wl_r<47> b_wl_r<46> b_wl_r<45> b_wl_r<44> b_wl_r<43> b_wl_r<42> b_wl_r<41> b_wl_r<40> b_wl_r<39> b_wl_r<38> b_wl_r<37> b_wl_r<36> b_wl_r<35> b_wl_r<34> b_wl_r<33> b_wl_r<32> b_wl_r<31> b_wl_r<30> b_wl_r<29> b_wl_r<28> b_wl_r<27> b_wl_r<26> b_wl_r<25> b_wl_r<24> b_wl_r<23> b_wl_r<22> b_wl_r<21> b_wl_r<20> b_wl_r<19> b_wl_r<18> b_wl_r<17> b_wl_r<16> b_wl_r<15> b_wl_r<14> b_wl_r<13> b_wl_r<12> b_wl_r<11> b_wl_r<10> b_wl_r<9> b_wl_r<8> b_wl_r<7> b_wl_r<6> b_wl_r<5> b_wl_r<4> b_wl_r<3> b_wl_r<2> b_wl_r<1> b_wl_r<0> VDDARRAY! VSS! / RM_IHPSG13_256x8_c2_2P_MATRIX_pcell_1
XRAM<0> a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0> b_blc_l<15> b_blc_l<14> b_blc_l<13> b_blc_l<12> b_blc_l<11> b_blc_l<10> b_blc_l<9> b_blc_l<8> b_blc_l<7> b_blc_l<6> b_blc_l<5> b_blc_l<4> b_blc_l<3> b_blc_l<2> b_blc_l<1> b_blc_l<0> b_blt_l<15> b_blt_l<14> b_blt_l<13> b_blt_l<12> b_blt_l<11> b_blt_l<10> b_blt_l<9> b_blt_l<8> b_blt_l<7> b_blt_l<6> b_blt_l<5> b_blt_l<4> b_blt_l<3> b_blt_l<2> b_blt_l<1> b_blt_l<0> b_wl_l<63> b_wl_l<62> b_wl_l<61> b_wl_l<60> b_wl_l<59> b_wl_l<58> b_wl_l<57> b_wl_l<56> b_wl_l<55> b_wl_l<54> b_wl_l<53> b_wl_l<52> b_wl_l<51> b_wl_l<50> b_wl_l<49> b_wl_l<48> b_wl_l<47> b_wl_l<46> b_wl_l<45> b_wl_l<44> b_wl_l<43> b_wl_l<42> b_wl_l<41> b_wl_l<40> b_wl_l<39> b_wl_l<38> b_wl_l<37> b_wl_l<36> b_wl_l<35> b_wl_l<34> b_wl_l<33> b_wl_l<32> b_wl_l<31> b_wl_l<30> b_wl_l<29> b_wl_l<28> b_wl_l<27> b_wl_l<26> b_wl_l<25> b_wl_l<24> b_wl_l<23> b_wl_l<22> b_wl_l<21> b_wl_l<20> b_wl_l<19> b_wl_l<18> b_wl_l<17> b_wl_l<16> b_wl_l<15> b_wl_l<14> b_wl_l<13> b_wl_l<12> b_wl_l<11> b_wl_l<10> b_wl_l<9> b_wl_l<8> b_wl_l<7> b_wl_l<6> b_wl_l<5> b_wl_l<4> b_wl_l<3> b_wl_l<2> b_wl_l<1> b_wl_l<0> VDDARRAY! VSS! / RM_IHPSG13_256x8_c2_2P_MATRIX_pcell_1


XB_COLDRV<1> b_addr_col<1> b_addr_col<0> b_addr_col_r<1> b_addr_col_r<0> b_addr_dec<7> b_addr_dec<6> b_addr_dec<5> b_addr_dec<4> b_addr_dec<3> b_addr_dec<2> b_addr_dec<1> b_addr_dec<0> b_addr_dec_r<7> b_addr_dec_r<6> b_addr_dec_r<5> b_addr_dec_r<4> b_addr_dec_r<3> b_addr_dec_r<2> b_addr_dec_r<1> b_addr_dec_r<0> b_dclk b_dclk_p_r<0> b_rclk b_rclk_p_r<0> b_wclk b_wclk_p_r<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13X8
XB_COLDRV<0> b_addr_col<1> b_addr_col<0> b_addr_col_l<1> b_addr_col_l<0> b_addr_dec<7> b_addr_dec<6> b_addr_dec<5> b_addr_dec<4> b_addr_dec<3> b_addr_dec<2> b_addr_dec<1> b_addr_dec<0> b_addr_dec_l<7> b_addr_dec_l<6> b_addr_dec_l<5> b_addr_dec_l<4> b_addr_dec_l<3> b_addr_dec_l<2> b_addr_dec_l<1> b_addr_dec_l<0> b_dclk b_dclk_p_l<0> b_rclk b_rclk_p_l<0> b_wclk b_wclk_p_l<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13X8
XA_COLDRV<1> a_addr_col<1> a_addr_col<0> a_addr_col_r<1> a_addr_col_r<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_r<7> a_addr_dec_r<6> a_addr_dec_r<5> a_addr_dec_r<4> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> a_dclk a_dclk_p_r<0> a_rclk a_rclk_p_r<0> a_wclk a_wclk_p_r<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13X8
XA_COLDRV<0> a_addr_col<1> a_addr_col<0> a_addr_col_l<1> a_addr_col_l<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_l<7> a_addr_dec_l<6> a_addr_dec_l<5> a_addr_dec_l<4> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> a_dclk a_dclk_p_l<0> a_rclk a_rclk_p_l<0> a_wclk a_wclk_p_l<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13X8


XB_WLDRV<7> b_wi<63> b_wi<62> b_wi<61> b_wi<60> b_wi<59> b_wi<58> b_wi<57> b_wi<56> b_wi<55> b_wi<54> b_wi<53> b_wi<52> b_wi<51> b_wi<50> b_wi<49> b_wi<48> b_wl_r<63> b_wl_r<62> b_wl_r<61> b_wl_r<60> b_wl_r<59> b_wl_r<58> b_wl_r<57> b_wl_r<56> b_wl_r<55> b_wl_r<54> b_wl_r<53> b_wl_r<52> b_wl_r<51> b_wl_r<50> b_wl_r<49> b_wl_r<48>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<6> b_wi<47> b_wi<46> b_wi<45> b_wi<44> b_wi<43> b_wi<42> b_wi<41> b_wi<40> b_wi<39> b_wi<38> b_wi<37> b_wi<36> b_wi<35> b_wi<34> b_wi<33> b_wi<32> b_wl_r<47> b_wl_r<46> b_wl_r<45> b_wl_r<44> b_wl_r<43> b_wl_r<42> b_wl_r<41> b_wl_r<40> b_wl_r<39> b_wl_r<38> b_wl_r<37> b_wl_r<36> b_wl_r<35> b_wl_r<34> b_wl_r<33> b_wl_r<32>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<5> b_wi<31> b_wi<30> b_wi<29> b_wi<28> b_wi<27> b_wi<26> b_wi<25> b_wi<24> b_wi<23> b_wi<22> b_wi<21> b_wi<20> b_wi<19> b_wi<18> b_wi<17> b_wi<16> b_wl_r<31> b_wl_r<30> b_wl_r<29> b_wl_r<28> b_wl_r<27> b_wl_r<26> b_wl_r<25> b_wl_r<24> b_wl_r<23> b_wl_r<22> b_wl_r<21> b_wl_r<20> b_wl_r<19> b_wl_r<18> b_wl_r<17> b_wl_r<16>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<4> b_wi<15> b_wi<14> b_wi<13> b_wi<12> b_wi<11> b_wi<10> b_wi<9> b_wi<8> b_wi<7> b_wi<6> b_wi<5> b_wi<4> b_wi<3> b_wi<2> b_wi<1> b_wi<0> b_wl_r<15> b_wl_r<14> b_wl_r<13> b_wl_r<12> b_wl_r<11> b_wl_r<10> b_wl_r<9> b_wl_r<8> b_wl_r<7> b_wl_r<6> b_wl_r<5> b_wl_r<4> b_wl_r<3> b_wl_r<2> b_wl_r<1> b_wl_r<0>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<3> b_wi<63> b_wi<62> b_wi<61> b_wi<60> b_wi<59> b_wi<58> b_wi<57> b_wi<56> b_wi<55> b_wi<54> b_wi<53> b_wi<52> b_wi<51> b_wi<50> b_wi<49> b_wi<48> b_wl_l<63> b_wl_l<62> b_wl_l<61> b_wl_l<60> b_wl_l<59> b_wl_l<58> b_wl_l<57> b_wl_l<56> b_wl_l<55> b_wl_l<54> b_wl_l<53> b_wl_l<52> b_wl_l<51> b_wl_l<50> b_wl_l<49> b_wl_l<48>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<2> b_wi<47> b_wi<46> b_wi<45> b_wi<44> b_wi<43> b_wi<42> b_wi<41> b_wi<40> b_wi<39> b_wi<38> b_wi<37> b_wi<36> b_wi<35> b_wi<34> b_wi<33> b_wi<32> b_wl_l<47> b_wl_l<46> b_wl_l<45> b_wl_l<44> b_wl_l<43> b_wl_l<42> b_wl_l<41> b_wl_l<40> b_wl_l<39> b_wl_l<38> b_wl_l<37> b_wl_l<36> b_wl_l<35> b_wl_l<34> b_wl_l<33> b_wl_l<32>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<1> b_wi<31> b_wi<30> b_wi<29> b_wi<28> b_wi<27> b_wi<26> b_wi<25> b_wi<24> b_wi<23> b_wi<22> b_wi<21> b_wi<20> b_wi<19> b_wi<18> b_wi<17> b_wi<16> b_wl_l<31> b_wl_l<30> b_wl_l<29> b_wl_l<28> b_wl_l<27> b_wl_l<26> b_wl_l<25> b_wl_l<24> b_wl_l<23> b_wl_l<22> b_wl_l<21> b_wl_l<20> b_wl_l<19> b_wl_l<18> b_wl_l<17> b_wl_l<16>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XB_WLDRV<0> b_wi<15> b_wi<14> b_wi<13> b_wi<12> b_wi<11> b_wi<10> b_wi<9> b_wi<8> b_wi<7> b_wi<6> b_wi<5> b_wi<4> b_wi<3> b_wi<2> b_wi<1> b_wi<0> b_wl_l<15> b_wl_l<14> b_wl_l<13> b_wl_l<12> b_wl_l<11> b_wl_l<10> b_wl_l<9> b_wl_l<8> b_wl_l<7> b_wl_l<6> b_wl_l<5> b_wl_l<4> b_wl_l<3> b_wl_l<2> b_wl_l<1> b_wl_l<0>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<7> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<6> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<5> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<4> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<3> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<2> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<1> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8
XA_WLDRV<0> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0>  VDD! VSS! / RM_IHPSG13_256x8_c2_2P_WLDRV16X8


XB_CTRL b_aclk_n B_BIST_CLK B_BIST_MEN B_BIST_EN B_BIST_REN B_BIST_WEN b_tiel B_CLK B_MEN b_dclk b_eclk b_pulse_h b_pulse_l b_pulse b_rclk B_REN b_cs b_wclk B_WEN VDD! VSS! / RM_IHPSG13_256x8_c2_2P_CTRL
XA_CTRL a_aclk_n A_BIST_CLK A_BIST_MEN A_BIST_EN A_BIST_REN A_BIST_WEN a_tiel A_CLK A_MEN a_dclk a_eclk a_pulse_h a_pulse_l a_pulse a_rclk A_REN a_cs a_wclk A_WEN VDD! VSS! / RM_IHPSG13_256x8_c2_2P_CTRL


XB_ROWDEC b_addr_row<5> b_addr_row<4> b_addr_row<3> b_addr_row<2> b_addr_row<1> b_addr_row<0> b_cs b_eclk b_wi<63> b_wi<62> b_wi<61> b_wi<60> b_wi<59> b_wi<58> b_wi<57> b_wi<56> b_wi<55> b_wi<54> b_wi<53> b_wi<52> b_wi<51> b_wi<50> b_wi<49> b_wi<48> b_wi<47> b_wi<46> b_wi<45> b_wi<44> b_wi<43> b_wi<42> b_wi<41> b_wi<40> b_wi<39> b_wi<38> b_wi<37> b_wi<36> b_wi<35> b_wi<34> b_wi<33> b_wi<32> b_wi<31> b_wi<30> b_wi<29> b_wi<28> b_wi<27> b_wi<26> b_wi<25> b_wi<24> b_wi<23> b_wi<22> b_wi<21> b_wi<20> b_wi<19> b_wi<18> b_wi<17> b_wi<16> b_wi<15> b_wi<14> b_wi<13> b_wi<12> b_wi<11> b_wi<10> b_wi<9> b_wi<8> b_wi<7> b_wi<6> b_wi<5> b_wi<4> b_wi<3> b_wi<2> b_wi<1> b_wi<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_ROWDEC6
XA_ROWDEC a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> a_cs a_eclk a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_ROWDEC6
XB_ROWREG b_aclk_n B_ADDR<7> B_ADDR<6> B_ADDR<5> B_ADDR<4> B_ADDR<3> B_ADDR<2> b_addr_row<5> b_addr_row<4> b_addr_row<3> b_addr_row<2> b_addr_row<1> b_addr_row<0> B_BIST_ADDR<7> B_BIST_ADDR<6> B_BIST_ADDR<5> B_BIST_ADDR<4> B_BIST_ADDR<3> B_BIST_ADDR<2> B_BIST_EN VDD! VSS!  / RM_IHPSG13_256x8_c2_2P_ROWREG6
XA_ROWREG a_aclk_n A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_EN VDD! VSS!  / RM_IHPSG13_256x8_c2_2P_ROWREG6
XB_COLDEC b_aclk_n B_ADDR<1> B_ADDR<0> b_addr_col<1> b_addr_col<0> b_addr_dec<7> b_addr_dec<6> b_addr_dec<5> b_addr_dec<4> b_addr_dec<3> b_addr_dec<2> b_addr_dec<1> b_addr_dec<0> B_BIST_ADDR<1> B_BIST_ADDR<0> B_BIST_EN VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDEC2
XA_COLDEC a_aclk_n A_ADDR<1> A_ADDR<0> a_addr_col<1> a_addr_col<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_EN VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDEC2


XB_DLYH b_pulse b_pulse_h VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_pcell_2
XB_DLYL b_pulse_x b_pulse_l VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_pcell_3
XA_DLYH a_pulse a_pulse_h VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_pcell_2
XA_DLYL a_pulse_x a_pulse_l VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_pcell_3
XB_DLYMUX b_pulse_h B_DLY b_pulse_x VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_MUX
XA_DLYMUX a_pulse_h A_DLY a_pulse_x VDD! VSS! / RM_IHPSG13_256x8_c2_2P_DLY_MUX

XCOLCTRL<7> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<7> A_BIST_DIN<7> A_BIST_EN a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> A_BM<7> a_dclk_n_r<3> a_dclk_n_r<4> a_dclk_p_r<3> a_dclk_p_r<4> A_DOUT<7> A_DIN<7> a_rclk_n_r<3> a_rclk_n_r<4> a_rclk_p_r<3> a_rclk_p_r<4> a_tieh<7> a_wclk_n_r<3> a_wclk_n_r<4> a_wclk_p_r<3> a_wclk_p_r<4> b_addr_dec_r<3> b_addr_dec_r<2> b_addr_dec_r<1> b_addr_dec_r<0> B_BIST_BM<7> B_BIST_DIN<7> B_BIST_EN b_blc_r<15> b_blc_r<14> b_blc_r<13> b_blc_r<12> b_blt_r<15> b_blt_r<14> b_blt_r<13> b_blt_r<12> B_BM<7> b_dclk_n_r<3> b_dclk_n_r<4> b_dclk_p_r<3> b_dclk_p_r<4> B_DOUT<7> B_DIN<7> b_rclk_n_r<3> b_rclk_n_r<4> b_rclk_p_r<3> b_rclk_p_r<4> b_tieh<7> b_wclk_n_r<3> b_wclk_n_r<4> b_wclk_p_r<3> b_wclk_p_r<4> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<6> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<6> A_BIST_DIN<6> A_BIST_EN a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> A_BM<6> a_dclk_n_r<2> a_dclk_n_r<3> a_dclk_p_r<2> a_dclk_p_r<3> A_DOUT<6> A_DIN<6> a_rclk_n_r<2> a_rclk_n_r<3> a_rclk_p_r<2> a_rclk_p_r<3> a_tieh<6> a_wclk_n_r<2> a_wclk_n_r<3> a_wclk_p_r<2> a_wclk_p_r<3> b_addr_dec_r<3> b_addr_dec_r<2> b_addr_dec_r<1> b_addr_dec_r<0> B_BIST_BM<6> B_BIST_DIN<6> B_BIST_EN b_blc_r<11> b_blc_r<10> b_blc_r<9> b_blc_r<8> b_blt_r<11> b_blt_r<10> b_blt_r<9> b_blt_r<8> B_BM<6> b_dclk_n_r<2> b_dclk_n_r<3> b_dclk_p_r<2> b_dclk_p_r<3> B_DOUT<6> B_DIN<6> b_rclk_n_r<2> b_rclk_n_r<3> b_rclk_p_r<2> b_rclk_p_r<3> b_tieh<6> b_wclk_n_r<2> b_wclk_n_r<3> b_wclk_p_r<2> b_wclk_p_r<3> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<5> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<5> A_BIST_DIN<5> A_BIST_EN a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> A_BM<5> a_dclk_n_r<1> a_dclk_n_r<2> a_dclk_p_r<1> a_dclk_p_r<2> A_DOUT<5> A_DIN<5> a_rclk_n_r<1> a_rclk_n_r<2> a_rclk_p_r<1> a_rclk_p_r<2> a_tieh<5> a_wclk_n_r<1> a_wclk_n_r<2> a_wclk_p_r<1> a_wclk_p_r<2> b_addr_dec_r<3> b_addr_dec_r<2> b_addr_dec_r<1> b_addr_dec_r<0> B_BIST_BM<5> B_BIST_DIN<5> B_BIST_EN b_blc_r<7> b_blc_r<6> b_blc_r<5> b_blc_r<4> b_blt_r<7> b_blt_r<6> b_blt_r<5> b_blt_r<4> B_BM<5> b_dclk_n_r<1> b_dclk_n_r<2> b_dclk_p_r<1> b_dclk_p_r<2> B_DOUT<5> B_DIN<5> b_rclk_n_r<1> b_rclk_n_r<2> b_rclk_p_r<1> b_rclk_p_r<2> b_tieh<5> b_wclk_n_r<1> b_wclk_n_r<2> b_wclk_p_r<1> b_wclk_p_r<2> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<4> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<4> A_BIST_DIN<4> A_BIST_EN a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> A_BM<4> a_dclk_n_r<0> a_dclk_n_r<1> a_dclk_p_r<0> a_dclk_p_r<1> A_DOUT<4> A_DIN<4> a_rclk_n_r<0> a_rclk_n_r<1> a_rclk_p_r<0> a_rclk_p_r<1> a_tieh<4> a_wclk_n_r<0> a_wclk_n_r<1> a_wclk_p_r<0> a_wclk_p_r<1> b_addr_dec_r<3> b_addr_dec_r<2> b_addr_dec_r<1> b_addr_dec_r<0> B_BIST_BM<4> B_BIST_DIN<4> B_BIST_EN b_blc_r<3> b_blc_r<2> b_blc_r<1> b_blc_r<0> b_blt_r<3> b_blt_r<2> b_blt_r<1> b_blt_r<0> B_BM<4> b_dclk_n_r<0> b_dclk_n_r<1> b_dclk_p_r<0> b_dclk_p_r<1> B_DOUT<4> B_DIN<4> b_rclk_n_r<0> b_rclk_n_r<1> b_rclk_p_r<0> b_rclk_p_r<1> b_tieh<4> b_wclk_n_r<0> b_wclk_n_r<1> b_wclk_p_r<0> b_wclk_p_r<1> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<3> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<0> A_BIST_DIN<0> A_BIST_EN a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> A_BM<0> a_dclk_n_l<3> a_dclk_n_l<4> a_dclk_p_l<3> a_dclk_p_l<4> A_DOUT<0> A_DIN<0> a_rclk_n_l<3> a_rclk_n_l<4> a_rclk_p_l<3> a_rclk_p_l<4> a_tieh<0> a_wclk_n_l<3> a_wclk_n_l<4> a_wclk_p_l<3> a_wclk_p_l<4> b_addr_dec_l<3> b_addr_dec_l<2> b_addr_dec_l<1> b_addr_dec_l<0> B_BIST_BM<0> B_BIST_DIN<0> B_BIST_EN b_blc_l<15> b_blc_l<14> b_blc_l<13> b_blc_l<12> b_blt_l<15> b_blt_l<14> b_blt_l<13> b_blt_l<12> B_BM<0> b_dclk_n_l<3> b_dclk_n_l<4> b_dclk_p_l<3> b_dclk_p_l<4> B_DOUT<0> B_DIN<0> b_rclk_n_l<3> b_rclk_n_l<4> b_rclk_p_l<3> b_rclk_p_l<4> b_tieh<0> b_wclk_n_l<3> b_wclk_n_l<4> b_wclk_p_l<3> b_wclk_p_l<4> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<2> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<1> A_BIST_DIN<1> A_BIST_EN a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> A_BM<1> a_dclk_n_l<2> a_dclk_n_l<3> a_dclk_p_l<2> a_dclk_p_l<3> A_DOUT<1> A_DIN<1> a_rclk_n_l<2> a_rclk_n_l<3> a_rclk_p_l<2> a_rclk_p_l<3> a_tieh<1> a_wclk_n_l<2> a_wclk_n_l<3> a_wclk_p_l<2> a_wclk_p_l<3> b_addr_dec_l<3> b_addr_dec_l<2> b_addr_dec_l<1> b_addr_dec_l<0> B_BIST_BM<1> B_BIST_DIN<1> B_BIST_EN b_blc_l<11> b_blc_l<10> b_blc_l<9> b_blc_l<8> b_blt_l<11> b_blt_l<10> b_blt_l<9> b_blt_l<8> B_BM<1> b_dclk_n_l<2> b_dclk_n_l<3> b_dclk_p_l<2> b_dclk_p_l<3> B_DOUT<1> B_DIN<1> b_rclk_n_l<2> b_rclk_n_l<3> b_rclk_p_l<2> b_rclk_p_l<3> b_tieh<1> b_wclk_n_l<2> b_wclk_n_l<3> b_wclk_p_l<2> b_wclk_p_l<3> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<1> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<2> A_BIST_DIN<2> A_BIST_EN a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> A_BM<2> a_dclk_n_l<1> a_dclk_n_l<2> a_dclk_p_l<1> a_dclk_p_l<2> A_DOUT<2> A_DIN<2> a_rclk_n_l<1> a_rclk_n_l<2> a_rclk_p_l<1> a_rclk_p_l<2> a_tieh<2> a_wclk_n_l<1> a_wclk_n_l<2> a_wclk_p_l<1> a_wclk_p_l<2> b_addr_dec_l<3> b_addr_dec_l<2> b_addr_dec_l<1> b_addr_dec_l<0> B_BIST_BM<2> B_BIST_DIN<2> B_BIST_EN b_blc_l<7> b_blc_l<6> b_blc_l<5> b_blc_l<4> b_blt_l<7> b_blt_l<6> b_blt_l<5> b_blt_l<4> B_BM<2> b_dclk_n_l<1> b_dclk_n_l<2> b_dclk_p_l<1> b_dclk_p_l<2> B_DOUT<2> B_DIN<2> b_rclk_n_l<1> b_rclk_n_l<2> b_rclk_p_l<1> b_rclk_p_l<2> b_tieh<2> b_wclk_n_l<1> b_wclk_n_l<2> b_wclk_p_l<1> b_wclk_p_l<2> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2
XCOLCTRL<0> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<3> A_BIST_DIN<3> A_BIST_EN a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> A_BM<3> a_dclk_n_l<0> a_dclk_n_l<1> a_dclk_p_l<0> a_dclk_p_l<1> A_DOUT<3> A_DIN<3> a_rclk_n_l<0> a_rclk_n_l<1> a_rclk_p_l<0> a_rclk_p_l<1> a_tieh<3> a_wclk_n_l<0> a_wclk_n_l<1> a_wclk_p_l<0> a_wclk_p_l<1> b_addr_dec_l<3> b_addr_dec_l<2> b_addr_dec_l<1> b_addr_dec_l<0> B_BIST_BM<3> B_BIST_DIN<3> B_BIST_EN b_blc_l<3> b_blc_l<2> b_blc_l<1> b_blc_l<0> b_blt_l<3> b_blt_l<2> b_blt_l<1> b_blt_l<0> B_BM<3> b_dclk_n_l<0> b_dclk_n_l<1> b_dclk_p_l<0> b_dclk_p_l<1> B_DOUT<3> B_DIN<3> b_rclk_n_l<0> b_rclk_n_l<1> b_rclk_p_l<0> b_rclk_p_l<1> b_tieh<3> b_wclk_n_l<0> b_wclk_n_l<1> b_wclk_p_l<0> b_wclk_p_l<1> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLCTRL2


XDRVFILL4<1> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<2> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<3> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<4> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<5> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<6> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<7> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<8> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<9> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XDRVFILL4<10> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4
XCOLFILL4<1> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<2> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<3> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<4> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<5> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<6> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<7> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<8> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<9> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<10> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<11> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<12> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<13> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<14> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<15> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<16> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<17> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<18> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<19> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<20> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<21> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<22> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<23> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
XCOLFILL4<24> VDD! VSS! / RM_IHPSG13_256x8_c2_2P_COLDRV13_FILL4C2
.ENDS
