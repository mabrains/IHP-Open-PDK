# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 13:36:37 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_256x8_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_256x8_c2_bm_bist 0 0 ;
  SIZE 278.51 BY 136.97 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.33 0 213.59 0.26 ;
    END
  END A_DIN[4]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.84 0 214.1 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 222 0 222.26 0.26 ;
    END
  END A_BM[4]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 220.625 0 220.885 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.19 0 206.45 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.88 0 216.14 0.26 ;
    END
  END B_DIN[4]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.35 0 214.61 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.365 0 207.625 0.26 ;
    END
  END B_BM[4]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 208.895 0 209.155 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.02 0 223.28 0.26 ;
    END
  END B_DOUT[4]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 259.105 0 263.525 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 241.425 0 245.845 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.745 0 228.165 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.065 0 210.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 176.475 0 179.285 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.175 0 168.985 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.725 0 153.535 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 140.425 0 143.235 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.275 0 138.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.975 0 127.785 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.525 0 112.335 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.225 0 102.035 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 136.97 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 267.945 0 272.365 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 250.265 0 254.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 232.585 0 237.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.905 0 219.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 171.325 0 174.135 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.025 0 163.835 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 155.875 0 158.685 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.575 0 148.385 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 130.125 0 132.935 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.825 0 122.635 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.675 0 117.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 104.375 0 107.185 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 267.945 53.41 272.365 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 250.265 53.41 254.685 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 232.585 53.41 237.005 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.905 53.41 219.325 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 136.97 ;
    END
  END VDDARRAY!
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.01 0 231.27 0.26 ;
    END
  END A_DIN[5]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.52 0 231.78 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 239.68 0 239.94 0.26 ;
    END
  END A_BM[5]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 238.305 0 238.565 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.87 0 224.13 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 233.56 0 233.82 0.26 ;
    END
  END B_DIN[5]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.03 0 232.29 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 225.045 0 225.305 0.26 ;
    END
  END B_BM[5]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.575 0 226.835 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 240.7 0 240.96 0.26 ;
    END
  END B_DOUT[5]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.69 0 248.95 0.26 ;
    END
  END A_DIN[6]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.2 0 249.46 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 257.36 0 257.62 0.26 ;
    END
  END A_BM[6]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 255.985 0 256.245 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.55 0 241.81 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 251.24 0 251.5 0.26 ;
    END
  END B_DIN[6]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.71 0 249.97 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 242.725 0 242.985 0.26 ;
    END
  END B_BM[6]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 244.255 0 244.515 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.38 0 258.64 0.26 ;
    END
  END B_DOUT[6]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.37 0 266.63 0.26 ;
    END
  END A_DIN[7]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.88 0 267.14 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 275.04 0 275.3 0.26 ;
    END
  END A_BM[7]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 273.665 0 273.925 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.23 0 259.49 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 268.92 0 269.18 0.26 ;
    END
  END B_DIN[7]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.39 0 267.65 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 260.405 0 260.665 0.26 ;
    END
  END B_BM[7]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 261.935 0 262.195 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.06 0 276.32 0.26 ;
    END
  END B_DOUT[7]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.345 0 155.605 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.955 0 161.215 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.905 0 123.165 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.295 0 117.555 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.855 0 156.115 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.465 0 161.725 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.395 0 122.655 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.785 0 117.045 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 164.525 0 164.785 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 165.035 0 165.295 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 113.725 0 113.985 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 113.215 0 113.475 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 163.505 0 163.765 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 164.015 0 164.275 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 114.745 0 115.005 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 114.235 0 114.495 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.125 0 144.385 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.635 0 144.895 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.125 0 134.385 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.615 0 133.875 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.105 0 143.365 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.615 0 143.875 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.145 0 135.405 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.635 0 134.895 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.075 0 167.335 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 166.565 0 166.825 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.175 0 111.435 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.685 0 111.945 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 166.055 0 166.315 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 165.545 0 165.805 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.195 0 112.455 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.705 0 112.965 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.815 0 154.075 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.385 0 157.645 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.875 0 157.135 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 154.325 0 154.585 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 174.725 0 174.985 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.435 0 124.695 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 120.865 0 121.125 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 121.375 0 121.635 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.925 0 124.185 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.525 0 103.785 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 96.5171 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.01 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.813443 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.365 0 156.625 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.285 0 152.545 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.915 0 159.175 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.405 0 158.665 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.795 0 153.055 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 97.0942 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.01 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.871096 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 121.885 0 122.145 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.965 0 126.225 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.335 0 119.595 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.845 0 120.105 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.455 0 125.715 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 278.51 136.97 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 136.94 ;
      RECT 1.135 136.21 1.335 136.94 ;
      RECT 1.545 136.21 1.905 136.94 ;
      RECT 2.115 136.21 2.315 136.94 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 136.21 2.97 136.94 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 136.21 3.54 136.94 ;
      RECT 3.835 136.21 4.035 136.94 ;
      RECT 4.33 136.21 4.69 136.94 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 136.21 5.1 136.94 ;
      RECT 5.555 136.21 5.755 136.94 ;
      RECT 5.965 136.21 6.325 136.94 ;
      RECT 6.535 136.21 6.735 136.94 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 136.21 7.39 136.94 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 136.21 7.96 136.94 ;
      RECT 8.255 136.21 8.455 136.94 ;
      RECT 8.75 136.21 9.11 136.94 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 136.21 9.52 136.94 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 136.21 10.175 136.94 ;
      RECT 10.385 136.21 10.745 136.94 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 136.21 11.155 136.94 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 136.21 11.81 136.94 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 136.21 12.38 136.94 ;
      RECT 12.675 136.21 12.875 136.94 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 136.21 13.53 136.94 ;
      RECT 13.74 136.21 13.94 136.94 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 136.21 14.595 136.94 ;
      RECT 14.805 136.21 15.165 136.94 ;
      RECT 15.375 136.21 15.575 136.94 ;
      RECT 16.03 136.21 16.23 136.94 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 136.21 16.8 136.94 ;
      RECT 17.095 136.21 17.295 136.94 ;
      RECT 17.59 136.21 17.95 136.94 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 136.21 18.36 136.94 ;
      RECT 18.815 136.21 19.015 136.94 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 136.21 19.585 136.94 ;
      RECT 19.795 136.21 19.995 136.94 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 136.21 20.65 136.94 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 136.21 21.22 136.94 ;
      RECT 21.515 136.21 21.715 136.94 ;
      RECT 22.01 136.21 22.37 136.94 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 136.21 22.78 136.94 ;
      RECT 23.235 136.21 23.435 136.94 ;
      RECT 23.645 136.21 24.005 136.94 ;
      RECT 24.215 136.21 24.415 136.94 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 136.21 25.07 136.94 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 136.21 25.64 136.94 ;
      RECT 25.935 136.21 26.135 136.94 ;
      RECT 26.43 136.21 26.79 136.94 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 136.21 27.2 136.94 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 136.21 27.855 136.94 ;
      RECT 28.065 136.21 28.425 136.94 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 136.21 28.835 136.94 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 136.21 29.49 136.94 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 136.21 30.06 136.94 ;
      RECT 30.355 136.21 30.555 136.94 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 136.21 31.21 136.94 ;
      RECT 31.42 136.21 31.62 136.94 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 136.21 32.275 136.94 ;
      RECT 32.485 136.21 32.845 136.94 ;
      RECT 33.055 136.21 33.255 136.94 ;
      RECT 33.71 136.21 33.91 136.94 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 136.21 34.48 136.94 ;
      RECT 34.775 136.21 34.975 136.94 ;
      RECT 35.27 136.21 35.63 136.94 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 136.21 36.04 136.94 ;
      RECT 36.495 136.21 36.695 136.94 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 136.21 37.265 136.94 ;
      RECT 37.475 136.21 37.675 136.94 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 136.21 38.33 136.94 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 136.21 38.9 136.94 ;
      RECT 39.195 136.21 39.395 136.94 ;
      RECT 39.69 136.21 40.05 136.94 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 136.21 40.46 136.94 ;
      RECT 40.915 136.21 41.115 136.94 ;
      RECT 41.325 136.21 41.685 136.94 ;
      RECT 41.895 136.21 42.095 136.94 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 136.21 42.75 136.94 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 136.21 43.32 136.94 ;
      RECT 43.615 136.21 43.815 136.94 ;
      RECT 44.11 136.21 44.47 136.94 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 136.21 44.88 136.94 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 136.21 45.535 136.94 ;
      RECT 45.745 136.21 46.105 136.94 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 136.21 46.515 136.94 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 136.21 47.17 136.94 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 136.21 47.74 136.94 ;
      RECT 48.035 136.21 48.235 136.94 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 136.21 48.89 136.94 ;
      RECT 49.1 136.21 49.3 136.94 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 136.21 49.955 136.94 ;
      RECT 50.165 136.21 50.525 136.94 ;
      RECT 50.735 136.21 50.935 136.94 ;
      RECT 51.39 136.21 51.59 136.94 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 136.21 52.16 136.94 ;
      RECT 52.455 136.21 52.655 136.94 ;
      RECT 52.95 136.21 53.31 136.94 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 136.21 53.72 136.94 ;
      RECT 54.175 136.21 54.375 136.94 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 136.21 54.945 136.94 ;
      RECT 55.155 136.21 55.355 136.94 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 136.21 56.01 136.94 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 136.21 56.58 136.94 ;
      RECT 56.875 136.21 57.075 136.94 ;
      RECT 57.37 136.21 57.73 136.94 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 136.21 58.14 136.94 ;
      RECT 58.595 136.21 58.795 136.94 ;
      RECT 59.005 136.21 59.365 136.94 ;
      RECT 59.575 136.21 59.775 136.94 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 136.21 60.43 136.94 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 136.21 61 136.94 ;
      RECT 61.295 136.21 61.495 136.94 ;
      RECT 61.79 136.21 62.15 136.94 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 136.21 62.56 136.94 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 136.21 63.215 136.94 ;
      RECT 63.425 136.21 63.785 136.94 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 136.21 64.195 136.94 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 136.21 64.85 136.94 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 136.21 65.42 136.94 ;
      RECT 65.715 136.21 65.915 136.94 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 136.21 66.57 136.94 ;
      RECT 66.78 136.21 66.98 136.94 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 136.21 67.635 136.94 ;
      RECT 67.845 136.21 68.205 136.94 ;
      RECT 68.415 136.21 68.615 136.94 ;
      RECT 69.07 136.21 69.27 136.94 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 136.21 69.84 136.94 ;
      RECT 70.135 136.21 70.335 136.94 ;
      RECT 70.63 136.21 70.99 136.94 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 136.21 71.4 136.94 ;
      RECT 71.855 136.21 72.055 136.94 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 73.59 0.17 74.36 0.43 ;
      RECT 73.59 0.17 73.85 8.7 ;
      RECT 74.1 0.17 74.36 8.7 ;
      RECT 74.61 0.18 75.38 0.88 ;
      RECT 74.61 0.18 74.87 8.7 ;
      RECT 75.12 0.18 75.38 8.7 ;
      RECT 75.63 0.17 76.4 0.43 ;
      RECT 75.63 0.17 75.89 8.7 ;
      RECT 76.14 0.17 76.4 8.7 ;
      RECT 76.65 0.18 77.42 0.88 ;
      RECT 76.65 0.18 76.91 8.7 ;
      RECT 77.16 0.18 77.42 8.7 ;
      RECT 77.67 0.17 78.44 0.43 ;
      RECT 77.67 0.17 77.93 8.7 ;
      RECT 78.18 0.17 78.44 8.7 ;
      RECT 78.69 0.18 79.46 0.88 ;
      RECT 78.69 0.18 78.95 8.7 ;
      RECT 79.2 0.18 79.46 8.7 ;
      RECT 79.71 0.17 80.48 0.43 ;
      RECT 79.71 0.17 79.97 8.7 ;
      RECT 80.22 0.17 80.48 8.7 ;
      RECT 80.73 0.18 81.5 0.88 ;
      RECT 80.73 0.18 80.99 8.7 ;
      RECT 81.24 0.18 81.5 8.7 ;
      RECT 81.75 0.17 82.52 0.43 ;
      RECT 81.75 0.17 82.01 8.7 ;
      RECT 82.26 0.17 82.52 8.7 ;
      RECT 82.77 0.18 83.54 0.88 ;
      RECT 82.77 0.18 83.03 8.7 ;
      RECT 83.28 0.18 83.54 8.7 ;
      RECT 83.79 0.17 84.56 0.43 ;
      RECT 83.79 0.17 84.05 8.7 ;
      RECT 84.3 0.17 84.56 8.7 ;
      RECT 84.81 0.18 85.58 0.88 ;
      RECT 84.81 0.18 85.07 8.7 ;
      RECT 85.32 0.18 85.58 8.7 ;
      RECT 85.83 0.17 86.6 0.43 ;
      RECT 85.83 0.17 86.09 8.7 ;
      RECT 86.34 0.17 86.6 8.7 ;
      RECT 86.85 0.18 87.62 0.88 ;
      RECT 86.85 0.18 87.11 8.7 ;
      RECT 87.36 0.18 87.62 8.7 ;
      RECT 87.87 0.17 88.64 0.43 ;
      RECT 87.87 0.17 88.13 8.7 ;
      RECT 88.38 0.17 88.64 8.7 ;
      RECT 88.89 0.18 89.66 0.88 ;
      RECT 88.89 0.18 89.15 8.7 ;
      RECT 89.4 0.18 89.66 8.7 ;
      RECT 89.91 0.17 90.68 0.43 ;
      RECT 89.91 0.17 90.17 8.7 ;
      RECT 90.42 0.17 90.68 8.7 ;
      RECT 90.93 0.18 91.7 0.88 ;
      RECT 90.93 0.18 91.19 8.7 ;
      RECT 91.44 0.18 91.7 8.7 ;
      RECT 91.95 0.17 92.72 0.43 ;
      RECT 91.95 0.17 92.21 8.7 ;
      RECT 92.46 0.17 92.72 8.7 ;
      RECT 92.97 0.18 93.74 0.88 ;
      RECT 92.97 0.18 93.23 8.7 ;
      RECT 93.48 0.18 93.74 8.7 ;
      RECT 93.99 0.17 94.76 0.43 ;
      RECT 93.99 0.17 94.25 8.7 ;
      RECT 94.5 0.17 94.76 8.7 ;
      RECT 95.01 0.18 95.78 0.88 ;
      RECT 95.01 0.18 95.27 8.7 ;
      RECT 95.52 0.18 95.78 8.7 ;
      RECT 96.03 0.17 96.8 0.43 ;
      RECT 96.03 0.17 96.29 8.7 ;
      RECT 96.54 0.17 96.8 8.7 ;
      RECT 97.05 0.18 97.82 0.88 ;
      RECT 97.05 0.18 97.31 8.7 ;
      RECT 97.56 0.18 97.82 8.7 ;
      RECT 72.265 136.21 72.625 136.94 ;
      RECT 72.835 136.21 73.035 136.94 ;
      RECT 99.445 0.18 100.215 0.88 ;
      RECT 99.445 0.18 99.705 8.7 ;
      RECT 99.955 0.18 100.215 8.7 ;
      RECT 100.465 0.17 101.235 0.43 ;
      RECT 100.465 0.17 100.725 8.7 ;
      RECT 100.975 0.17 101.235 8.7 ;
      RECT 73.66 136.13 73.86 136.94 ;
      RECT 98.425 0.3 98.685 8.7 ;
      RECT 102.505 0.18 103.275 0.88 ;
      RECT 102.505 0.18 102.765 8.7 ;
      RECT 103.015 0.18 103.275 8.7 ;
      RECT 98.935 0.3 99.195 8.7 ;
      RECT 101.485 0 101.745 8.7 ;
      RECT 101.995 0 102.255 8.7 ;
      RECT 103.525 0.52 103.785 8.7 ;
      RECT 104.035 0.3 104.295 8.7 ;
      RECT 104.545 0.3 104.805 8.7 ;
      RECT 105.055 0.3 105.315 8.7 ;
      RECT 105.565 0.3 105.825 8.7 ;
      RECT 106.075 0.3 106.335 8.7 ;
      RECT 106.585 0.3 106.845 8.7 ;
      RECT 107.095 0.3 107.355 8.7 ;
      RECT 109.135 0.18 109.905 0.88 ;
      RECT 109.135 0.18 109.395 8.7 ;
      RECT 109.645 0.18 109.905 8.7 ;
      RECT 107.605 0.3 107.865 8.7 ;
      RECT 108.115 0 108.375 8.7 ;
      RECT 108.625 0 108.885 8.7 ;
      RECT 110.155 0 110.415 8.7 ;
      RECT 110.665 0 110.925 8.7 ;
      RECT 111.175 0.52 111.435 8.7 ;
      RECT 111.685 0.52 111.945 8.7 ;
      RECT 112.195 0.52 112.455 8.7 ;
      RECT 112.705 0.52 112.965 8.7 ;
      RECT 113.215 0.52 113.475 8.7 ;
      RECT 113.725 0.52 113.985 8.7 ;
      RECT 114.235 0.52 114.495 8.7 ;
      RECT 114.745 0.52 115.005 8.7 ;
      RECT 115.255 0.3 115.515 8.7 ;
      RECT 115.765 0.3 116.025 8.7 ;
      RECT 116.275 0.3 116.535 8.7 ;
      RECT 116.785 0.52 117.045 8.7 ;
      RECT 117.295 0.52 117.555 8.7 ;
      RECT 117.805 0.3 118.065 8.7 ;
      RECT 118.315 0.3 118.575 8.7 ;
      RECT 118.825 0.3 119.085 8.7 ;
      RECT 119.335 0.52 119.595 8.7 ;
      RECT 119.845 0.52 120.105 8.7 ;
      RECT 120.355 0.3 120.615 8.7 ;
      RECT 120.865 0.52 121.125 8.7 ;
      RECT 121.375 0.52 121.635 8.7 ;
      RECT 121.885 0.52 122.145 8.7 ;
      RECT 122.395 0.52 122.655 8.7 ;
      RECT 122.905 0.52 123.165 8.7 ;
      RECT 123.415 0.3 123.675 8.7 ;
      RECT 123.925 0.52 124.185 8.7 ;
      RECT 124.435 0.52 124.695 8.7 ;
      RECT 124.945 0.3 125.205 8.7 ;
      RECT 125.455 0.52 125.715 8.7 ;
      RECT 127.495 0.17 128.265 0.43 ;
      RECT 127.495 0.17 127.755 8.7 ;
      RECT 128.005 0.17 128.265 8.7 ;
      RECT 125.965 0.52 126.225 8.7 ;
      RECT 126.475 0.3 126.735 8.7 ;
      RECT 126.985 0.3 127.245 8.7 ;
      RECT 130.045 0.17 130.815 0.43 ;
      RECT 130.045 0.17 130.305 8.7 ;
      RECT 130.555 0.17 130.815 8.7 ;
      RECT 128.515 0.3 128.775 8.7 ;
      RECT 131.575 0.18 132.345 0.88 ;
      RECT 131.575 0.18 131.835 8.7 ;
      RECT 132.085 0.18 132.345 8.7 ;
      RECT 129.025 0.3 129.285 8.7 ;
      RECT 129.535 0.3 129.795 8.7 ;
      RECT 131.065 0.3 131.325 8.7 ;
      RECT 132.595 0 132.855 8.7 ;
      RECT 133.105 0 133.365 8.7 ;
      RECT 133.615 0.52 133.875 8.7 ;
      RECT 134.125 0.52 134.385 8.7 ;
      RECT 134.635 0.52 134.895 8.7 ;
      RECT 135.145 0.52 135.405 8.7 ;
      RECT 135.655 0 135.915 8.7 ;
      RECT 136.165 0 136.425 8.7 ;
      RECT 136.675 0.3 136.935 8.7 ;
      RECT 137.185 0.3 137.445 8.7 ;
      RECT 137.695 0 137.955 8.7 ;
      RECT 138.205 0 138.465 8.7 ;
      RECT 138.715 0.3 138.975 8.7 ;
      RECT 139.535 0.3 139.795 8.7 ;
      RECT 140.045 0 140.305 8.7 ;
      RECT 140.555 0 140.815 8.7 ;
      RECT 141.065 0.3 141.325 8.7 ;
      RECT 141.575 0.3 141.835 8.7 ;
      RECT 142.085 0 142.345 8.7 ;
      RECT 142.595 0 142.855 8.7 ;
      RECT 143.105 0.52 143.365 8.7 ;
      RECT 143.615 0.52 143.875 8.7 ;
      RECT 144.125 0.52 144.385 8.7 ;
      RECT 146.165 0.18 146.935 0.88 ;
      RECT 146.165 0.18 146.425 8.7 ;
      RECT 146.675 0.18 146.935 8.7 ;
      RECT 144.635 0.52 144.895 8.7 ;
      RECT 147.695 0.17 148.465 0.43 ;
      RECT 147.695 0.17 147.955 8.7 ;
      RECT 148.205 0.17 148.465 8.7 ;
      RECT 145.145 0 145.405 8.7 ;
      RECT 145.655 0 145.915 8.7 ;
      RECT 147.185 0.3 147.445 8.7 ;
      RECT 150.245 0.17 151.015 0.43 ;
      RECT 150.245 0.17 150.505 8.7 ;
      RECT 150.755 0.17 151.015 8.7 ;
      RECT 148.715 0.3 148.975 8.7 ;
      RECT 149.225 0.3 149.485 8.7 ;
      RECT 149.735 0.3 149.995 8.7 ;
      RECT 151.265 0.3 151.525 8.7 ;
      RECT 151.775 0.3 152.035 8.7 ;
      RECT 152.285 0.52 152.545 8.7 ;
      RECT 152.795 0.52 153.055 8.7 ;
      RECT 153.305 0.3 153.565 8.7 ;
      RECT 153.815 0.52 154.075 8.7 ;
      RECT 154.325 0.52 154.585 8.7 ;
      RECT 154.835 0.3 155.095 8.7 ;
      RECT 155.345 0.52 155.605 8.7 ;
      RECT 155.855 0.52 156.115 8.7 ;
      RECT 156.365 0.52 156.625 8.7 ;
      RECT 156.875 0.52 157.135 8.7 ;
      RECT 157.385 0.52 157.645 8.7 ;
      RECT 157.895 0.3 158.155 8.7 ;
      RECT 158.405 0.52 158.665 8.7 ;
      RECT 158.915 0.52 159.175 8.7 ;
      RECT 159.425 0.3 159.685 8.7 ;
      RECT 159.935 0.3 160.195 8.7 ;
      RECT 160.445 0.3 160.705 8.7 ;
      RECT 160.955 0.52 161.215 8.7 ;
      RECT 161.465 0.52 161.725 8.7 ;
      RECT 161.975 0.3 162.235 8.7 ;
      RECT 162.485 0.3 162.745 8.7 ;
      RECT 162.995 0.3 163.255 8.7 ;
      RECT 163.505 0.52 163.765 8.7 ;
      RECT 164.015 0.52 164.275 8.7 ;
      RECT 164.525 0.52 164.785 8.7 ;
      RECT 165.035 0.52 165.295 8.7 ;
      RECT 165.545 0.52 165.805 8.7 ;
      RECT 166.055 0.52 166.315 8.7 ;
      RECT 166.565 0.52 166.825 8.7 ;
      RECT 168.605 0.18 169.375 0.88 ;
      RECT 168.605 0.18 168.865 8.7 ;
      RECT 169.115 0.18 169.375 8.7 ;
      RECT 167.075 0.52 167.335 8.7 ;
      RECT 167.585 0 167.845 8.7 ;
      RECT 168.095 0 168.355 8.7 ;
      RECT 169.625 0 169.885 8.7 ;
      RECT 170.135 0 170.395 8.7 ;
      RECT 170.645 0.3 170.905 8.7 ;
      RECT 171.155 0.3 171.415 8.7 ;
      RECT 171.665 0.3 171.925 8.7 ;
      RECT 172.175 0.3 172.435 8.7 ;
      RECT 172.685 0.3 172.945 8.7 ;
      RECT 173.195 0.3 173.455 8.7 ;
      RECT 175.235 0.18 176.005 0.88 ;
      RECT 175.235 0.18 175.495 8.7 ;
      RECT 175.745 0.18 176.005 8.7 ;
      RECT 173.705 0.3 173.965 8.7 ;
      RECT 174.215 0.3 174.475 8.7 ;
      RECT 177.275 0.17 178.045 0.43 ;
      RECT 177.275 0.17 177.535 8.7 ;
      RECT 177.785 0.17 178.045 8.7 ;
      RECT 178.295 0.18 179.065 0.88 ;
      RECT 178.295 0.18 178.555 8.7 ;
      RECT 178.805 0.18 179.065 8.7 ;
      RECT 174.725 0.52 174.985 8.7 ;
      RECT 176.255 0 176.515 8.7 ;
      RECT 180.69 0.18 181.46 0.88 ;
      RECT 180.69 0.18 180.95 8.7 ;
      RECT 181.2 0.18 181.46 8.7 ;
      RECT 181.71 0.17 182.48 0.43 ;
      RECT 181.71 0.17 181.97 8.7 ;
      RECT 182.22 0.17 182.48 8.7 ;
      RECT 182.73 0.18 183.5 0.88 ;
      RECT 182.73 0.18 182.99 8.7 ;
      RECT 183.24 0.18 183.5 8.7 ;
      RECT 183.75 0.17 184.52 0.43 ;
      RECT 183.75 0.17 184.01 8.7 ;
      RECT 184.26 0.17 184.52 8.7 ;
      RECT 184.77 0.18 185.54 0.88 ;
      RECT 184.77 0.18 185.03 8.7 ;
      RECT 185.28 0.18 185.54 8.7 ;
      RECT 185.79 0.17 186.56 0.43 ;
      RECT 185.79 0.17 186.05 8.7 ;
      RECT 186.3 0.17 186.56 8.7 ;
      RECT 186.81 0.18 187.58 0.88 ;
      RECT 186.81 0.18 187.07 8.7 ;
      RECT 187.32 0.18 187.58 8.7 ;
      RECT 187.83 0.17 188.6 0.43 ;
      RECT 187.83 0.17 188.09 8.7 ;
      RECT 188.34 0.17 188.6 8.7 ;
      RECT 188.85 0.18 189.62 0.88 ;
      RECT 188.85 0.18 189.11 8.7 ;
      RECT 189.36 0.18 189.62 8.7 ;
      RECT 189.87 0.17 190.64 0.43 ;
      RECT 189.87 0.17 190.13 8.7 ;
      RECT 190.38 0.17 190.64 8.7 ;
      RECT 190.89 0.18 191.66 0.88 ;
      RECT 190.89 0.18 191.15 8.7 ;
      RECT 191.4 0.18 191.66 8.7 ;
      RECT 191.91 0.17 192.68 0.43 ;
      RECT 191.91 0.17 192.17 8.7 ;
      RECT 192.42 0.17 192.68 8.7 ;
      RECT 192.93 0.18 193.7 0.88 ;
      RECT 192.93 0.18 193.19 8.7 ;
      RECT 193.44 0.18 193.7 8.7 ;
      RECT 193.95 0.17 194.72 0.43 ;
      RECT 193.95 0.17 194.21 8.7 ;
      RECT 194.46 0.17 194.72 8.7 ;
      RECT 194.97 0.18 195.74 0.88 ;
      RECT 194.97 0.18 195.23 8.7 ;
      RECT 195.48 0.18 195.74 8.7 ;
      RECT 195.99 0.17 196.76 0.43 ;
      RECT 195.99 0.17 196.25 8.7 ;
      RECT 196.5 0.17 196.76 8.7 ;
      RECT 197.01 0.18 197.78 0.88 ;
      RECT 197.01 0.18 197.27 8.7 ;
      RECT 197.52 0.18 197.78 8.7 ;
      RECT 198.03 0.17 198.8 0.43 ;
      RECT 198.03 0.17 198.29 8.7 ;
      RECT 198.54 0.17 198.8 8.7 ;
      RECT 199.05 0.18 199.82 0.88 ;
      RECT 199.05 0.18 199.31 8.7 ;
      RECT 199.56 0.18 199.82 8.7 ;
      RECT 200.07 0.17 200.84 0.43 ;
      RECT 200.07 0.17 200.33 8.7 ;
      RECT 200.58 0.17 200.84 8.7 ;
      RECT 201.09 0.18 201.86 0.88 ;
      RECT 201.09 0.18 201.35 8.7 ;
      RECT 201.6 0.18 201.86 8.7 ;
      RECT 202.11 0.17 202.88 0.43 ;
      RECT 202.11 0.17 202.37 8.7 ;
      RECT 202.62 0.17 202.88 8.7 ;
      RECT 203.13 0.18 203.9 0.88 ;
      RECT 203.13 0.18 203.39 8.7 ;
      RECT 203.64 0.18 203.9 8.7 ;
      RECT 176.765 0 177.025 8.7 ;
      RECT 204.15 0.17 204.92 0.43 ;
      RECT 204.15 0.17 204.41 8.7 ;
      RECT 204.66 0.17 204.92 8.7 ;
      RECT 179.315 0.3 179.575 8.7 ;
      RECT 179.825 0.3 180.085 8.7 ;
      RECT 204.65 136.13 204.85 136.94 ;
      RECT 205.475 136.21 205.675 136.94 ;
      RECT 205.885 136.21 206.245 136.94 ;
      RECT 206.19 0.52 206.45 4.315 ;
      RECT 206.455 136.21 206.655 136.94 ;
      RECT 207.11 136.21 207.31 136.94 ;
      RECT 207.365 0.52 207.625 2.82 ;
      RECT 207.52 136.21 207.88 136.94 ;
      RECT 208.175 136.21 208.375 136.94 ;
      RECT 208.67 136.21 209.03 136.94 ;
      RECT 209.605 0.18 210.375 0.88 ;
      RECT 209.605 0.18 209.865 12.9 ;
      RECT 210.115 0.18 210.375 12.9 ;
      RECT 208.895 0.52 209.155 2.82 ;
      RECT 209.24 136.21 209.44 136.94 ;
      RECT 210.625 0.155 211.395 0.445 ;
      RECT 210.625 0.155 210.885 13.21 ;
      RECT 211.135 0.155 211.395 13.21 ;
      RECT 209.895 136.21 210.095 136.94 ;
      RECT 210.305 136.21 210.665 136.94 ;
      RECT 210.875 136.21 211.075 136.94 ;
      RECT 211.53 136.21 211.73 136.94 ;
      RECT 211.94 136.21 212.3 136.94 ;
      RECT 212.595 136.21 212.795 136.94 ;
      RECT 213.09 136.21 213.45 136.94 ;
      RECT 213.33 0.52 213.59 14.115 ;
      RECT 213.66 136.21 213.86 136.94 ;
      RECT 213.84 0.52 214.1 13.45 ;
      RECT 214.315 136.21 214.515 136.94 ;
      RECT 214.86 0.155 215.63 0.445 ;
      RECT 214.86 0.155 215.12 8.665 ;
      RECT 215.37 0.155 215.63 8.665 ;
      RECT 214.35 0.52 214.61 11.315 ;
      RECT 214.725 136.21 215.085 136.94 ;
      RECT 215.295 136.21 215.495 136.94 ;
      RECT 215.88 0.52 216.14 9.955 ;
      RECT 215.95 136.21 216.15 136.94 ;
      RECT 216.36 136.21 216.72 136.94 ;
      RECT 217.015 136.21 217.215 136.94 ;
      RECT 217.51 136.21 217.87 136.94 ;
      RECT 217.92 0.3 218.18 8.7 ;
      RECT 218.08 136.21 218.28 136.94 ;
      RECT 218.735 136.21 218.935 136.94 ;
      RECT 218.43 0.18 219.2 0.88 ;
      RECT 219.145 136.21 219.505 136.94 ;
      RECT 219.715 136.21 219.915 136.94 ;
      RECT 220.37 136.21 220.57 136.94 ;
      RECT 220.625 0.52 220.885 6.28 ;
      RECT 220.78 136.21 221.14 136.94 ;
      RECT 221.435 136.21 221.635 136.94 ;
      RECT 222 0.52 222.26 5.57 ;
      RECT 221.93 136.21 222.29 136.94 ;
      RECT 222.5 136.21 222.7 136.94 ;
      RECT 222.51 0.3 222.77 5.235 ;
      RECT 223.02 0.52 223.28 7.78 ;
      RECT 223.155 136.21 223.355 136.94 ;
      RECT 223.565 136.21 223.925 136.94 ;
      RECT 223.87 0.52 224.13 4.315 ;
      RECT 224.135 136.21 224.335 136.94 ;
      RECT 224.79 136.21 224.99 136.94 ;
      RECT 225.045 0.52 225.305 2.82 ;
      RECT 225.2 136.21 225.56 136.94 ;
      RECT 225.855 136.21 226.055 136.94 ;
      RECT 226.35 136.21 226.71 136.94 ;
      RECT 227.285 0.18 228.055 0.88 ;
      RECT 227.285 0.18 227.545 12.9 ;
      RECT 227.795 0.18 228.055 12.9 ;
      RECT 226.575 0.52 226.835 2.82 ;
      RECT 226.92 136.21 227.12 136.94 ;
      RECT 228.305 0.155 229.075 0.445 ;
      RECT 228.305 0.155 228.565 13.21 ;
      RECT 228.815 0.155 229.075 13.21 ;
      RECT 227.575 136.21 227.775 136.94 ;
      RECT 227.985 136.21 228.345 136.94 ;
      RECT 228.555 136.21 228.755 136.94 ;
      RECT 229.21 136.21 229.41 136.94 ;
      RECT 229.62 136.21 229.98 136.94 ;
      RECT 230.275 136.21 230.475 136.94 ;
      RECT 230.77 136.21 231.13 136.94 ;
      RECT 231.01 0.52 231.27 14.115 ;
      RECT 231.34 136.21 231.54 136.94 ;
      RECT 231.52 0.52 231.78 13.45 ;
      RECT 231.995 136.21 232.195 136.94 ;
      RECT 232.54 0.155 233.31 0.445 ;
      RECT 232.54 0.155 232.8 8.665 ;
      RECT 233.05 0.155 233.31 8.665 ;
      RECT 232.03 0.52 232.29 11.315 ;
      RECT 232.405 136.21 232.765 136.94 ;
      RECT 232.975 136.21 233.175 136.94 ;
      RECT 233.56 0.52 233.82 9.955 ;
      RECT 233.63 136.21 233.83 136.94 ;
      RECT 234.04 136.21 234.4 136.94 ;
      RECT 234.695 136.21 234.895 136.94 ;
      RECT 235.19 136.21 235.55 136.94 ;
      RECT 235.6 0.3 235.86 8.7 ;
      RECT 235.76 136.21 235.96 136.94 ;
      RECT 236.415 136.21 236.615 136.94 ;
      RECT 236.11 0.18 236.88 0.88 ;
      RECT 236.825 136.21 237.185 136.94 ;
      RECT 237.395 136.21 237.595 136.94 ;
      RECT 238.05 136.21 238.25 136.94 ;
      RECT 238.305 0.52 238.565 6.28 ;
      RECT 238.46 136.21 238.82 136.94 ;
      RECT 239.115 136.21 239.315 136.94 ;
      RECT 239.68 0.52 239.94 5.57 ;
      RECT 239.61 136.21 239.97 136.94 ;
      RECT 240.18 136.21 240.38 136.94 ;
      RECT 240.19 0.3 240.45 5.235 ;
      RECT 240.7 0.52 240.96 7.78 ;
      RECT 240.835 136.21 241.035 136.94 ;
      RECT 241.245 136.21 241.605 136.94 ;
      RECT 241.55 0.52 241.81 4.315 ;
      RECT 241.815 136.21 242.015 136.94 ;
      RECT 242.47 136.21 242.67 136.94 ;
      RECT 242.725 0.52 242.985 2.82 ;
      RECT 242.88 136.21 243.24 136.94 ;
      RECT 243.535 136.21 243.735 136.94 ;
      RECT 244.03 136.21 244.39 136.94 ;
      RECT 244.965 0.18 245.735 0.88 ;
      RECT 244.965 0.18 245.225 12.9 ;
      RECT 245.475 0.18 245.735 12.9 ;
      RECT 244.255 0.52 244.515 2.82 ;
      RECT 244.6 136.21 244.8 136.94 ;
      RECT 245.985 0.155 246.755 0.445 ;
      RECT 245.985 0.155 246.245 13.21 ;
      RECT 246.495 0.155 246.755 13.21 ;
      RECT 245.255 136.21 245.455 136.94 ;
      RECT 245.665 136.21 246.025 136.94 ;
      RECT 246.235 136.21 246.435 136.94 ;
      RECT 246.89 136.21 247.09 136.94 ;
      RECT 247.3 136.21 247.66 136.94 ;
      RECT 247.955 136.21 248.155 136.94 ;
      RECT 248.45 136.21 248.81 136.94 ;
      RECT 248.69 0.52 248.95 14.115 ;
      RECT 249.02 136.21 249.22 136.94 ;
      RECT 249.2 0.52 249.46 13.45 ;
      RECT 249.675 136.21 249.875 136.94 ;
      RECT 250.22 0.155 250.99 0.445 ;
      RECT 250.22 0.155 250.48 8.665 ;
      RECT 250.73 0.155 250.99 8.665 ;
      RECT 249.71 0.52 249.97 11.315 ;
      RECT 250.085 136.21 250.445 136.94 ;
      RECT 250.655 136.21 250.855 136.94 ;
      RECT 251.24 0.52 251.5 9.955 ;
      RECT 251.31 136.21 251.51 136.94 ;
      RECT 251.72 136.21 252.08 136.94 ;
      RECT 252.375 136.21 252.575 136.94 ;
      RECT 252.87 136.21 253.23 136.94 ;
      RECT 253.28 0.3 253.54 8.7 ;
      RECT 253.44 136.21 253.64 136.94 ;
      RECT 254.095 136.21 254.295 136.94 ;
      RECT 253.79 0.18 254.56 0.88 ;
      RECT 254.505 136.21 254.865 136.94 ;
      RECT 255.075 136.21 255.275 136.94 ;
      RECT 255.73 136.21 255.93 136.94 ;
      RECT 255.985 0.52 256.245 6.28 ;
      RECT 256.14 136.21 256.5 136.94 ;
      RECT 256.795 136.21 256.995 136.94 ;
      RECT 257.36 0.52 257.62 5.57 ;
      RECT 257.29 136.21 257.65 136.94 ;
      RECT 257.86 136.21 258.06 136.94 ;
      RECT 257.87 0.3 258.13 5.235 ;
      RECT 258.38 0.52 258.64 7.78 ;
      RECT 258.515 136.21 258.715 136.94 ;
      RECT 258.925 136.21 259.285 136.94 ;
      RECT 259.23 0.52 259.49 4.315 ;
      RECT 259.495 136.21 259.695 136.94 ;
      RECT 260.15 136.21 260.35 136.94 ;
      RECT 260.405 0.52 260.665 2.82 ;
      RECT 260.56 136.21 260.92 136.94 ;
      RECT 261.215 136.21 261.415 136.94 ;
      RECT 261.71 136.21 262.07 136.94 ;
      RECT 262.645 0.18 263.415 0.88 ;
      RECT 262.645 0.18 262.905 12.9 ;
      RECT 263.155 0.18 263.415 12.9 ;
      RECT 261.935 0.52 262.195 2.82 ;
      RECT 262.28 136.21 262.48 136.94 ;
      RECT 263.665 0.155 264.435 0.445 ;
      RECT 263.665 0.155 263.925 13.21 ;
      RECT 264.175 0.155 264.435 13.21 ;
      RECT 262.935 136.21 263.135 136.94 ;
      RECT 263.345 136.21 263.705 136.94 ;
      RECT 263.915 136.21 264.115 136.94 ;
      RECT 264.57 136.21 264.77 136.94 ;
      RECT 264.98 136.21 265.34 136.94 ;
      RECT 265.635 136.21 265.835 136.94 ;
      RECT 266.13 136.21 266.49 136.94 ;
      RECT 266.37 0.52 266.63 14.115 ;
      RECT 266.7 136.21 266.9 136.94 ;
      RECT 266.88 0.52 267.14 13.45 ;
      RECT 267.355 136.21 267.555 136.94 ;
      RECT 267.9 0.155 268.67 0.445 ;
      RECT 267.9 0.155 268.16 8.665 ;
      RECT 268.41 0.155 268.67 8.665 ;
      RECT 267.39 0.52 267.65 11.315 ;
      RECT 267.765 136.21 268.125 136.94 ;
      RECT 268.335 136.21 268.535 136.94 ;
      RECT 268.92 0.52 269.18 9.955 ;
      RECT 268.99 136.21 269.19 136.94 ;
      RECT 269.4 136.21 269.76 136.94 ;
      RECT 270.055 136.21 270.255 136.94 ;
      RECT 270.55 136.21 270.91 136.94 ;
      RECT 270.96 0.3 271.22 8.7 ;
      RECT 271.12 136.21 271.32 136.94 ;
      RECT 271.775 136.21 271.975 136.94 ;
      RECT 271.47 0.18 272.24 0.88 ;
      RECT 272.185 136.21 272.545 136.94 ;
      RECT 272.755 136.21 272.955 136.94 ;
      RECT 273.41 136.21 273.61 136.94 ;
      RECT 273.665 0.52 273.925 6.28 ;
      RECT 273.82 136.21 274.18 136.94 ;
      RECT 274.475 136.21 274.675 136.94 ;
      RECT 275.04 0.52 275.3 5.57 ;
      RECT 274.97 136.21 275.33 136.94 ;
      RECT 275.54 136.21 275.74 136.94 ;
      RECT 275.55 0.3 275.81 5.235 ;
      RECT 276.06 0.52 276.32 7.78 ;
      RECT 276.195 136.21 276.395 136.94 ;
      RECT 276.605 136.21 276.965 136.94 ;
      RECT 277.175 136.21 277.375 136.94 ;
      RECT 278 53.41 278.2 136.94 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 274.185 0 274.78 136.97 ;
      RECT 275.55 0.3 275.81 136.97 ;
      RECT 276.58 0 278.51 136.97 ;
      RECT 0 0.52 278.51 136.97 ;
      RECT 269.44 0 273.405 136.97 ;
      RECT 267.9 0.155 268.67 136.97 ;
      RECT 262.455 0 266.11 136.97 ;
      RECT 260.925 0 261.675 136.97 ;
      RECT 259.75 0 260.145 136.97 ;
      RECT 257.87 0.3 258.13 136.97 ;
      RECT 256.505 0 257.1 136.97 ;
      RECT 251.76 0 255.725 136.97 ;
      RECT 250.22 0.155 250.99 136.97 ;
      RECT 244.775 0 248.43 136.97 ;
      RECT 243.245 0 243.995 136.97 ;
      RECT 242.07 0 242.465 136.97 ;
      RECT 240.19 0.3 240.45 136.97 ;
      RECT 238.825 0 239.42 136.97 ;
      RECT 234.08 0 238.045 136.97 ;
      RECT 232.54 0.155 233.31 136.97 ;
      RECT 227.095 0 230.75 136.97 ;
      RECT 225.565 0 226.315 136.97 ;
      RECT 224.39 0 224.785 136.97 ;
      RECT 222.51 0.3 222.77 136.97 ;
      RECT 221.145 0 221.74 136.97 ;
      RECT 216.4 0 220.365 136.97 ;
      RECT 214.86 0.155 215.63 136.97 ;
      RECT 209.415 0 213.07 136.97 ;
      RECT 207.885 0 208.635 136.97 ;
      RECT 206.71 0 207.105 136.97 ;
      RECT 175.235 0.18 205.93 136.97 ;
      RECT 175.245 0 205.93 136.97 ;
      RECT 167.585 0.3 174.475 136.97 ;
      RECT 161.975 0.3 163.255 136.97 ;
      RECT 159.425 0.3 160.705 136.97 ;
      RECT 157.895 0.3 158.155 136.97 ;
      RECT 154.835 0.3 155.095 136.97 ;
      RECT 153.305 0.3 153.565 136.97 ;
      RECT 145.145 0.3 152.035 136.97 ;
      RECT 135.655 0 142.855 136.97 ;
      RECT 126.475 0.3 133.365 136.97 ;
      RECT 126.485 0 133.365 136.97 ;
      RECT 124.945 0.3 125.205 136.97 ;
      RECT 123.415 0.3 123.675 136.97 ;
      RECT 120.355 0.3 120.615 136.97 ;
      RECT 117.805 0.3 119.085 136.97 ;
      RECT 115.255 0.3 116.535 136.97 ;
      RECT 104.035 0.3 110.925 136.97 ;
      RECT 104.045 0 110.925 136.97 ;
      RECT 72.58 0.18 103.275 136.97 ;
      RECT 71.405 0 71.8 136.97 ;
      RECT 69.875 0 70.625 136.97 ;
      RECT 65.44 0 69.095 136.97 ;
      RECT 62.88 0.155 63.65 136.97 ;
      RECT 58.145 0 62.11 136.97 ;
      RECT 56.77 0 57.365 136.97 ;
      RECT 55.74 0.3 56 136.97 ;
      RECT 53.725 0 54.12 136.97 ;
      RECT 52.195 0 52.945 136.97 ;
      RECT 47.76 0 51.415 136.97 ;
      RECT 45.2 0.155 45.97 136.97 ;
      RECT 40.465 0 44.43 136.97 ;
      RECT 39.09 0 39.685 136.97 ;
      RECT 38.06 0.3 38.32 136.97 ;
      RECT 36.045 0 36.44 136.97 ;
      RECT 34.515 0 35.265 136.97 ;
      RECT 30.08 0 33.735 136.97 ;
      RECT 27.52 0.155 28.29 136.97 ;
      RECT 22.785 0 26.75 136.97 ;
      RECT 21.41 0 22.005 136.97 ;
      RECT 20.38 0.3 20.64 136.97 ;
      RECT 18.365 0 18.76 136.97 ;
      RECT 16.835 0 17.585 136.97 ;
      RECT 12.4 0 16.055 136.97 ;
      RECT 9.84 0.155 10.61 136.97 ;
      RECT 5.105 0 9.07 136.97 ;
      RECT 3.73 0 4.325 136.97 ;
      RECT 2.7 0.3 2.96 136.97 ;
      RECT 0 0 1.93 136.97 ;
      RECT 275.56 0 275.8 136.97 ;
      RECT 257.88 0 258.12 136.97 ;
      RECT 240.2 0 240.44 136.97 ;
      RECT 222.52 0 222.76 136.97 ;
      RECT 167.585 0 174.465 136.97 ;
      RECT 161.985 0 163.245 136.97 ;
      RECT 159.435 0 160.695 136.97 ;
      RECT 157.905 0 158.145 136.97 ;
      RECT 154.845 0 155.085 136.97 ;
      RECT 153.315 0 153.555 136.97 ;
      RECT 145.145 0 152.025 136.97 ;
      RECT 124.955 0 125.195 136.97 ;
      RECT 123.425 0 123.665 136.97 ;
      RECT 120.365 0 120.605 136.97 ;
      RECT 117.815 0 119.075 136.97 ;
      RECT 115.265 0 116.525 136.97 ;
      RECT 55.75 0 55.99 136.97 ;
      RECT 38.07 0 38.31 136.97 ;
      RECT 20.39 0 20.63 136.97 ;
      RECT 2.71 0 2.95 136.97 ;
      RECT 72.58 0 103.265 136.97 ;
      RECT 267.91 0 268.66 136.97 ;
      RECT 250.23 0 250.98 136.97 ;
      RECT 232.55 0 233.3 136.97 ;
      RECT 214.87 0 215.62 136.97 ;
      RECT 62.89 0 63.64 136.97 ;
      RECT 45.21 0 45.96 136.97 ;
      RECT 27.53 0 28.28 136.97 ;
      RECT 9.85 0 10.6 136.97 ;
    LAYER Metal3 ;
      RECT 0 0 278.51 136.97 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 179.545 0 205.805 136.97 ;
      RECT 174.395 0 176.215 136.97 ;
      RECT 169.245 0 171.065 136.97 ;
      RECT 272.625 0 278.51 136.97 ;
      RECT 263.785 0 267.685 136.97 ;
      RECT 263.785 47.305 278.51 53.15 ;
      RECT 254.945 0 258.845 136.97 ;
      RECT 246.105 0 250.005 136.97 ;
      RECT 246.105 47.305 258.845 53.15 ;
      RECT 237.265 0 241.165 136.97 ;
      RECT 228.425 0 232.325 136.97 ;
      RECT 228.425 47.305 241.165 53.15 ;
      RECT 219.585 0 223.485 136.97 ;
      RECT 210.745 0 214.645 136.97 ;
      RECT 210.745 47.305 223.485 53.15 ;
      RECT 164.095 0 165.915 136.97 ;
      RECT 158.945 0 160.765 136.97 ;
      RECT 153.795 0 155.615 136.97 ;
      RECT 148.645 0 150.465 136.97 ;
      RECT 143.495 0 145.315 136.97 ;
      RECT 138.345 0 140.165 136.97 ;
      RECT 133.195 0 135.015 136.97 ;
      RECT 128.045 0 129.865 136.97 ;
      RECT 122.895 0 124.715 136.97 ;
      RECT 117.745 0 119.565 136.97 ;
      RECT 112.595 0 114.415 136.97 ;
      RECT 107.445 0 109.265 136.97 ;
      RECT 102.295 0 104.115 136.97 ;
      RECT 72.705 0 98.965 136.97 ;
      RECT 63.865 0 67.765 136.97 ;
      RECT 55.025 0 58.925 136.97 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 136.97 ;
      RECT 37.345 0 41.245 136.97 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 136.97 ;
      RECT 19.665 0 23.565 136.97 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 136.97 ;
      RECT 0 0 5.885 136.97 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_256x8_c2_bm_bist

END LIBRARY
