# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 13:09:02 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_1024x32_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_1024x32_c2_bm_bist 0 0 ;
  SIZE 685.49 BY 385.37 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 408.15 0 408.41 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.08 0 277.34 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 408.66 0 408.92 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.57 0 276.83 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 416.82 0 417.08 0.26 ;
    END
  END A_BM[16]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 268.41 0 268.67 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 415.445 0 415.705 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 269.785 0 270.045 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.01 0 401.27 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.22 0 284.48 0.26 ;
    END
  END A_DOUT[15]
  PIN B_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 410.7 0 410.96 0.26 ;
    END
  END B_DIN[16]
  PIN B_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 274.53 0 274.79 0.26 ;
    END
  END B_DIN[15]
  PIN B_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 409.17 0 409.43 0.26 ;
    END
  END B_BIST_DIN[16]
  PIN B_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.06 0 276.32 0.26 ;
    END
  END B_BIST_DIN[15]
  PIN B_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 402.185 0 402.445 0.26 ;
    END
  END B_BM[16]
  PIN B_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 283.045 0 283.305 0.26 ;
    END
  END B_BM[15]
  PIN B_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 403.715 0 403.975 0.26 ;
    END
  END B_BIST_BM[16]
  PIN B_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 281.515 0 281.775 0.26 ;
    END
  END B_BIST_BM[15]
  PIN B_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 417.84 0 418.1 0.26 ;
    END
  END B_DOUT[16]
  PIN B_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.39 0 267.65 0.26 ;
    END
  END B_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 666.085 0 670.505 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.405 0 652.825 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 630.725 0 635.145 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 613.045 0 617.465 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.365 0 599.785 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 577.685 0 582.105 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.005 0 564.425 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 542.325 0 546.745 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.645 0 529.065 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.965 0 511.385 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 489.285 0 493.705 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 471.605 0 476.025 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 453.925 0 458.345 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 436.245 0 440.665 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 418.565 0 422.985 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 400.885 0 405.305 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 379.965 0 382.775 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.665 0 372.475 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.215 0 357.025 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 343.915 0 346.725 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 338.765 0 341.575 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 328.465 0 331.275 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.015 0 315.825 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.715 0 305.525 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.185 0 284.605 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.505 0 266.925 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 244.825 0 249.245 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 227.145 0 231.565 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.465 0 213.885 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 191.785 0 196.205 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.105 0 178.525 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.425 0 160.845 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.745 0 143.165 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.065 0 125.485 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.385 0 107.805 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.705 0 90.125 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 385.37 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 674.925 0 679.345 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 657.245 0 661.665 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.565 0 643.985 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.885 0 626.305 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 604.205 0 608.625 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.525 0 590.945 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.845 0 573.265 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 551.165 0 555.585 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.485 0 537.905 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.805 0 520.225 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 498.125 0 502.545 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.445 0 484.865 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.765 0 467.185 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 445.085 0 449.505 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.405 0 431.825 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.725 0 414.145 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 374.815 0 377.625 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.515 0 367.325 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 359.365 0 362.175 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 349.065 0 351.875 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.615 0 336.425 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 323.315 0 326.125 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 318.165 0 320.975 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 307.865 0 310.675 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 0 275.765 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 0 258.085 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 0 240.405 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 0 222.725 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 0 205.045 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 0 187.365 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 0 169.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 0 152.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 0 134.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 0 116.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 0 98.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 0 81.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 674.925 53.41 679.345 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 657.245 53.41 661.665 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.565 53.41 643.985 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.885 53.41 626.305 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 604.205 53.41 608.625 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.525 53.41 590.945 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.845 53.41 573.265 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 551.165 53.41 555.585 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.485 53.41 537.905 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.805 53.41 520.225 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 498.125 53.41 502.545 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.445 53.41 484.865 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.765 53.41 467.185 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 445.085 53.41 449.505 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.405 53.41 431.825 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.725 53.41 414.145 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 53.41 275.765 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 53.41 258.085 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 53.41 240.405 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 53.41 222.725 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 53.41 205.045 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 53.41 187.365 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 53.41 169.685 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 53.41 152.005 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 53.41 134.325 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 53.41 116.645 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 53.41 98.965 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 53.41 81.285 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 385.37 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 385.37 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 425.83 0 426.09 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.4 0 259.66 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 426.34 0 426.6 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.89 0 259.15 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 434.5 0 434.76 0.26 ;
    END
  END A_BM[17]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 250.73 0 250.99 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 433.125 0 433.385 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 252.105 0 252.365 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 418.69 0 418.95 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.54 0 266.8 0.26 ;
    END
  END A_DOUT[14]
  PIN B_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 428.38 0 428.64 0.26 ;
    END
  END B_DIN[17]
  PIN B_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 256.85 0 257.11 0.26 ;
    END
  END B_DIN[14]
  PIN B_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 426.85 0 427.11 0.26 ;
    END
  END B_BIST_DIN[17]
  PIN B_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.38 0 258.64 0.26 ;
    END
  END B_BIST_DIN[14]
  PIN B_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 419.865 0 420.125 0.26 ;
    END
  END B_BM[17]
  PIN B_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 265.365 0 265.625 0.26 ;
    END
  END B_BM[14]
  PIN B_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 421.395 0 421.655 0.26 ;
    END
  END B_BIST_BM[17]
  PIN B_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 263.835 0 264.095 0.26 ;
    END
  END B_BIST_BM[14]
  PIN B_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 435.52 0 435.78 0.26 ;
    END
  END B_DOUT[17]
  PIN B_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.71 0 249.97 0.26 ;
    END
  END B_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 443.51 0 443.77 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.72 0 241.98 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 444.02 0 444.28 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.21 0 241.47 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 452.18 0 452.44 0.26 ;
    END
  END A_BM[18]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 233.05 0 233.31 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 450.805 0 451.065 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 234.425 0 234.685 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 436.37 0 436.63 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.86 0 249.12 0.26 ;
    END
  END A_DOUT[13]
  PIN B_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 446.06 0 446.32 0.26 ;
    END
  END B_DIN[18]
  PIN B_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 239.17 0 239.43 0.26 ;
    END
  END B_DIN[13]
  PIN B_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 444.53 0 444.79 0.26 ;
    END
  END B_BIST_DIN[18]
  PIN B_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 240.7 0 240.96 0.26 ;
    END
  END B_BIST_DIN[13]
  PIN B_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 437.545 0 437.805 0.26 ;
    END
  END B_BM[18]
  PIN B_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 247.685 0 247.945 0.26 ;
    END
  END B_BM[13]
  PIN B_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 439.075 0 439.335 0.26 ;
    END
  END B_BIST_BM[18]
  PIN B_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 246.155 0 246.415 0.26 ;
    END
  END B_BIST_BM[13]
  PIN B_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 453.2 0 453.46 0.26 ;
    END
  END B_DOUT[18]
  PIN B_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.03 0 232.29 0.26 ;
    END
  END B_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.19 0 461.45 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.04 0 224.3 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.7 0 461.96 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.53 0 223.79 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 469.86 0 470.12 0.26 ;
    END
  END A_BM[19]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.37 0 215.63 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 468.485 0 468.745 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 216.745 0 217.005 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 454.05 0 454.31 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.18 0 231.44 0.26 ;
    END
  END A_DOUT[12]
  PIN B_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 463.74 0 464 0.26 ;
    END
  END B_DIN[19]
  PIN B_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221.49 0 221.75 0.26 ;
    END
  END B_DIN[12]
  PIN B_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 462.21 0 462.47 0.26 ;
    END
  END B_BIST_DIN[19]
  PIN B_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.02 0 223.28 0.26 ;
    END
  END B_BIST_DIN[12]
  PIN B_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 455.225 0 455.485 0.26 ;
    END
  END B_BM[19]
  PIN B_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 230.005 0 230.265 0.26 ;
    END
  END B_BM[12]
  PIN B_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 456.755 0 457.015 0.26 ;
    END
  END B_BIST_BM[19]
  PIN B_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.475 0 228.735 0.26 ;
    END
  END B_BIST_BM[12]
  PIN B_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 470.88 0 471.14 0.26 ;
    END
  END B_DOUT[19]
  PIN B_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.35 0 214.61 0.26 ;
    END
  END B_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 478.87 0 479.13 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.36 0 206.62 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 479.38 0 479.64 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.85 0 206.11 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 487.54 0 487.8 0.26 ;
    END
  END A_BM[20]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 197.69 0 197.95 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 486.165 0 486.425 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 199.065 0 199.325 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 471.73 0 471.99 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.5 0 213.76 0.26 ;
    END
  END A_DOUT[11]
  PIN B_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 481.42 0 481.68 0.26 ;
    END
  END B_DIN[20]
  PIN B_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.81 0 204.07 0.26 ;
    END
  END B_DIN[11]
  PIN B_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 479.89 0 480.15 0.26 ;
    END
  END B_BIST_DIN[20]
  PIN B_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.34 0 205.6 0.26 ;
    END
  END B_BIST_DIN[11]
  PIN B_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 472.905 0 473.165 0.26 ;
    END
  END B_BM[20]
  PIN B_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 212.325 0 212.585 0.26 ;
    END
  END B_BM[11]
  PIN B_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 474.435 0 474.695 0.26 ;
    END
  END B_BIST_BM[20]
  PIN B_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 210.795 0 211.055 0.26 ;
    END
  END B_BIST_BM[11]
  PIN B_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 488.56 0 488.82 0.26 ;
    END
  END B_DOUT[20]
  PIN B_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.67 0 196.93 0.26 ;
    END
  END B_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 496.55 0 496.81 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.68 0 188.94 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 497.06 0 497.32 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.17 0 188.43 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 505.22 0 505.48 0.26 ;
    END
  END A_BM[21]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 180.01 0 180.27 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 503.845 0 504.105 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.385 0 181.645 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 489.41 0 489.67 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.82 0 196.08 0.26 ;
    END
  END A_DOUT[10]
  PIN B_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 499.1 0 499.36 0.26 ;
    END
  END B_DIN[21]
  PIN B_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 186.13 0 186.39 0.26 ;
    END
  END B_DIN[10]
  PIN B_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 497.57 0 497.83 0.26 ;
    END
  END B_BIST_DIN[21]
  PIN B_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 187.66 0 187.92 0.26 ;
    END
  END B_BIST_DIN[10]
  PIN B_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 490.585 0 490.845 0.26 ;
    END
  END B_BM[21]
  PIN B_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 194.645 0 194.905 0.26 ;
    END
  END B_BM[10]
  PIN B_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 492.115 0 492.375 0.26 ;
    END
  END B_BIST_BM[21]
  PIN B_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.115 0 193.375 0.26 ;
    END
  END B_BIST_BM[10]
  PIN B_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 506.24 0 506.5 0.26 ;
    END
  END B_DOUT[21]
  PIN B_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.99 0 179.25 0.26 ;
    END
  END B_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.23 0 514.49 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171 0 171.26 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.74 0 515 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 170.49 0 170.75 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 522.9 0 523.16 0.26 ;
    END
  END A_BM[22]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 162.33 0 162.59 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 521.525 0 521.785 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 163.705 0 163.965 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 507.09 0 507.35 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.14 0 178.4 0.26 ;
    END
  END A_DOUT[9]
  PIN B_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 516.78 0 517.04 0.26 ;
    END
  END B_DIN[22]
  PIN B_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.45 0 168.71 0.26 ;
    END
  END B_DIN[9]
  PIN B_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 515.25 0 515.51 0.26 ;
    END
  END B_BIST_DIN[22]
  PIN B_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 169.98 0 170.24 0.26 ;
    END
  END B_BIST_DIN[9]
  PIN B_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 508.265 0 508.525 0.26 ;
    END
  END B_BM[22]
  PIN B_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.965 0 177.225 0.26 ;
    END
  END B_BM[9]
  PIN B_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 509.795 0 510.055 0.26 ;
    END
  END B_BIST_BM[22]
  PIN B_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 175.435 0 175.695 0.26 ;
    END
  END B_BIST_BM[9]
  PIN B_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 523.92 0 524.18 0.26 ;
    END
  END B_DOUT[22]
  PIN B_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.31 0 161.57 0.26 ;
    END
  END B_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 531.91 0 532.17 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.32 0 153.58 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 532.42 0 532.68 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.81 0 153.07 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 540.58 0 540.84 0.26 ;
    END
  END A_BM[23]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.65 0 144.91 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 539.205 0 539.465 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.025 0 146.285 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 524.77 0 525.03 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.46 0 160.72 0.26 ;
    END
  END A_DOUT[8]
  PIN B_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 534.46 0 534.72 0.26 ;
    END
  END B_DIN[23]
  PIN B_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.77 0 151.03 0.26 ;
    END
  END B_DIN[8]
  PIN B_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 532.93 0 533.19 0.26 ;
    END
  END B_BIST_DIN[23]
  PIN B_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.3 0 152.56 0.26 ;
    END
  END B_BIST_DIN[8]
  PIN B_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 525.945 0 526.205 0.26 ;
    END
  END B_BM[23]
  PIN B_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 159.285 0 159.545 0.26 ;
    END
  END B_BM[8]
  PIN B_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 527.475 0 527.735 0.26 ;
    END
  END B_BIST_BM[23]
  PIN B_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.755 0 158.015 0.26 ;
    END
  END B_BIST_BM[8]
  PIN B_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 541.6 0 541.86 0.26 ;
    END
  END B_DOUT[23]
  PIN B_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.63 0 143.89 0.26 ;
    END
  END B_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 549.59 0 549.85 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.64 0 135.9 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 550.1 0 550.36 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.13 0 135.39 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 558.26 0 558.52 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.97 0 127.23 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 556.885 0 557.145 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 128.345 0 128.605 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 542.45 0 542.71 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.78 0 143.04 0.26 ;
    END
  END A_DOUT[7]
  PIN B_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 552.14 0 552.4 0.26 ;
    END
  END B_DIN[24]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.09 0 133.35 0.26 ;
    END
  END B_DIN[7]
  PIN B_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 550.61 0 550.87 0.26 ;
    END
  END B_BIST_DIN[24]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.62 0 134.88 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 543.625 0 543.885 0.26 ;
    END
  END B_BM[24]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 141.605 0 141.865 0.26 ;
    END
  END B_BM[7]
  PIN B_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 545.155 0 545.415 0.26 ;
    END
  END B_BIST_BM[24]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 140.075 0 140.335 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 559.28 0 559.54 0.26 ;
    END
  END B_DOUT[24]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.95 0 126.21 0.26 ;
    END
  END B_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 567.27 0 567.53 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.96 0 118.22 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 567.78 0 568.04 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.45 0 117.71 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 575.94 0 576.2 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.29 0 109.55 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 574.565 0 574.825 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.665 0 110.925 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 560.13 0 560.39 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.1 0 125.36 0.26 ;
    END
  END A_DOUT[6]
  PIN B_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 569.82 0 570.08 0.26 ;
    END
  END B_DIN[25]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.41 0 115.67 0.26 ;
    END
  END B_DIN[6]
  PIN B_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 568.29 0 568.55 0.26 ;
    END
  END B_BIST_DIN[25]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.94 0 117.2 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 561.305 0 561.565 0.26 ;
    END
  END B_BM[25]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.925 0 124.185 0.26 ;
    END
  END B_BM[6]
  PIN B_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 562.835 0 563.095 0.26 ;
    END
  END B_BIST_BM[25]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.395 0 122.655 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 576.96 0 577.22 0.26 ;
    END
  END B_DOUT[25]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.27 0 108.53 0.26 ;
    END
  END B_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 584.95 0 585.21 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.28 0 100.54 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.46 0 585.72 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.77 0 100.03 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 593.62 0 593.88 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 91.61 0 91.87 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 592.245 0 592.505 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 92.985 0 93.245 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 577.81 0 578.07 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 107.42 0 107.68 0.26 ;
    END
  END A_DOUT[5]
  PIN B_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 587.5 0 587.76 0.26 ;
    END
  END B_DIN[26]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 97.73 0 97.99 0.26 ;
    END
  END B_DIN[5]
  PIN B_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.97 0 586.23 0.26 ;
    END
  END B_BIST_DIN[26]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.26 0 99.52 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 578.985 0 579.245 0.26 ;
    END
  END B_BM[26]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 106.245 0 106.505 0.26 ;
    END
  END B_BM[5]
  PIN B_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 580.515 0 580.775 0.26 ;
    END
  END B_BIST_BM[26]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.715 0 104.975 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 594.64 0 594.9 0.26 ;
    END
  END B_DOUT[26]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 90.59 0 90.85 0.26 ;
    END
  END B_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 602.63 0 602.89 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.6 0 82.86 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 603.14 0 603.4 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.09 0 82.35 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 611.3 0 611.56 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 73.93 0 74.19 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 609.925 0 610.185 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 75.305 0 75.565 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 595.49 0 595.75 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.74 0 90 0.26 ;
    END
  END A_DOUT[4]
  PIN B_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 605.18 0 605.44 0.26 ;
    END
  END B_DIN[27]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 80.05 0 80.31 0.26 ;
    END
  END B_DIN[4]
  PIN B_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 603.65 0 603.91 0.26 ;
    END
  END B_BIST_DIN[27]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.58 0 81.84 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 596.665 0 596.925 0.26 ;
    END
  END B_BM[27]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.565 0 88.825 0.26 ;
    END
  END B_BM[4]
  PIN B_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 598.195 0 598.455 0.26 ;
    END
  END B_BIST_BM[27]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 87.035 0 87.295 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 612.32 0 612.58 0.26 ;
    END
  END B_DOUT[27]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.91 0 73.17 0.26 ;
    END
  END B_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 620.31 0 620.57 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 620.82 0 621.08 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 628.98 0 629.24 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 627.605 0 627.865 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 613.17 0 613.43 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 622.86 0 623.12 0.26 ;
    END
  END B_DIN[28]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 621.33 0 621.59 0.26 ;
    END
  END B_BIST_DIN[28]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 614.345 0 614.605 0.26 ;
    END
  END B_BM[28]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 615.875 0 616.135 0.26 ;
    END
  END B_BIST_BM[28]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 630 0 630.26 0.26 ;
    END
  END B_DOUT[28]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 637.99 0 638.25 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 638.5 0 638.76 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 646.66 0 646.92 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 645.285 0 645.545 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 630.85 0 631.11 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 640.54 0 640.8 0.26 ;
    END
  END B_DIN[29]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 639.01 0 639.27 0.26 ;
    END
  END B_BIST_DIN[29]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 632.025 0 632.285 0.26 ;
    END
  END B_BM[29]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 633.555 0 633.815 0.26 ;
    END
  END B_BIST_BM[29]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 647.68 0 647.94 0.26 ;
    END
  END B_DOUT[29]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 655.67 0 655.93 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 656.18 0 656.44 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 664.34 0 664.6 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 662.965 0 663.225 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 648.53 0 648.79 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 658.22 0 658.48 0.26 ;
    END
  END B_DIN[30]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 656.69 0 656.95 0.26 ;
    END
  END B_BIST_DIN[30]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 649.705 0 649.965 0.26 ;
    END
  END B_BM[30]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 651.235 0 651.495 0.26 ;
    END
  END B_BIST_BM[30]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 665.36 0 665.62 0.26 ;
    END
  END B_DOUT[30]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 673.35 0 673.61 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 673.86 0 674.12 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 682.02 0 682.28 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 680.645 0 680.905 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 666.21 0 666.47 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 675.9 0 676.16 0.26 ;
    END
  END B_DIN[31]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 674.37 0 674.63 0.26 ;
    END
  END B_BIST_DIN[31]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 667.385 0 667.645 0.26 ;
    END
  END B_BM[31]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 668.915 0 669.175 0.26 ;
    END
  END B_BIST_BM[31]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 683.04 0 683.3 0.26 ;
    END
  END B_DOUT[31]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 358.835 0 359.095 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.445 0 364.705 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 326.395 0 326.655 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 320.785 0 321.045 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 359.345 0 359.605 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.955 0 365.215 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 325.885 0 326.145 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 320.275 0 320.535 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 368.015 0 368.275 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 368.525 0 368.785 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 317.215 0 317.475 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 316.705 0 316.965 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 366.995 0 367.255 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 367.505 0 367.765 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 318.235 0 318.495 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 317.725 0 317.985 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.615 0 347.875 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 348.125 0 348.385 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.615 0 337.875 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.105 0 337.365 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.595 0 346.855 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.105 0 347.365 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.635 0 338.895 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.125 0 338.385 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 370.565 0 370.825 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 370.055 0 370.315 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 314.665 0 314.925 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.175 0 315.435 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.545 0 369.805 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.035 0 369.295 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.685 0 315.945 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 316.195 0 316.455 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.115 0 373.375 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.625 0 373.885 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN B_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 312.115 0 312.375 0.26 ;
    END
  END B_ADDR[8]
  PIN B_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.605 0 311.865 0.26 ;
    END
  END B_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.075 0 371.335 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.585 0 371.845 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN B_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 314.155 0 314.415 0.26 ;
    END
  END B_ADDR[9]
  PIN B_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7995 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 69.61165 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 313.645 0 313.905 0.26 ;
    END
  END B_BIST_ADDR[9]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 357.305 0 357.565 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.875 0 361.135 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.365 0 360.625 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 357.815 0 358.075 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.215 0 378.475 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.925 0 328.185 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 324.355 0 324.615 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 324.865 0 325.125 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.415 0 327.675 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 307.015 0 307.275 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 254.5589 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.885 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.300258 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 359.855 0 360.115 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.775 0 356.035 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.405 0 362.665 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 361.895 0 362.155 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.285 0 356.545 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 254.9981 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.885 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.316009 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 325.375 0 325.635 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 329.455 0 329.715 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 322.825 0 323.085 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 323.335 0 323.595 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 328.945 0 329.205 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 685.49 385.37 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 385.34 ;
      RECT 1.135 384.61 1.335 385.34 ;
      RECT 1.545 384.61 1.905 385.34 ;
      RECT 2.115 384.61 2.315 385.34 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 384.61 2.97 385.34 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 384.61 3.54 385.34 ;
      RECT 3.835 384.61 4.035 385.34 ;
      RECT 4.33 384.61 4.69 385.34 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 384.61 5.1 385.34 ;
      RECT 5.555 384.61 5.755 385.34 ;
      RECT 5.965 384.61 6.325 385.34 ;
      RECT 6.535 384.61 6.735 385.34 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 384.61 7.39 385.34 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 384.61 7.96 385.34 ;
      RECT 8.255 384.61 8.455 385.34 ;
      RECT 8.75 384.61 9.11 385.34 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 384.61 9.52 385.34 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 384.61 10.175 385.34 ;
      RECT 10.385 384.61 10.745 385.34 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 384.61 11.155 385.34 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 384.61 11.81 385.34 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 384.61 12.38 385.34 ;
      RECT 12.675 384.61 12.875 385.34 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 384.61 13.53 385.34 ;
      RECT 13.74 384.61 13.94 385.34 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 384.61 14.595 385.34 ;
      RECT 14.805 384.61 15.165 385.34 ;
      RECT 15.375 384.61 15.575 385.34 ;
      RECT 16.03 384.61 16.23 385.34 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 384.61 16.8 385.34 ;
      RECT 17.095 384.61 17.295 385.34 ;
      RECT 17.59 384.61 17.95 385.34 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 384.61 18.36 385.34 ;
      RECT 18.815 384.61 19.015 385.34 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 384.61 19.585 385.34 ;
      RECT 19.795 384.61 19.995 385.34 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 384.61 20.65 385.34 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 384.61 21.22 385.34 ;
      RECT 21.515 384.61 21.715 385.34 ;
      RECT 22.01 384.61 22.37 385.34 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 384.61 22.78 385.34 ;
      RECT 23.235 384.61 23.435 385.34 ;
      RECT 23.645 384.61 24.005 385.34 ;
      RECT 24.215 384.61 24.415 385.34 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 384.61 25.07 385.34 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 384.61 25.64 385.34 ;
      RECT 25.935 384.61 26.135 385.34 ;
      RECT 26.43 384.61 26.79 385.34 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 384.61 27.2 385.34 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 384.61 27.855 385.34 ;
      RECT 28.065 384.61 28.425 385.34 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 384.61 28.835 385.34 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 384.61 29.49 385.34 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 384.61 30.06 385.34 ;
      RECT 30.355 384.61 30.555 385.34 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 384.61 31.21 385.34 ;
      RECT 31.42 384.61 31.62 385.34 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 384.61 32.275 385.34 ;
      RECT 32.485 384.61 32.845 385.34 ;
      RECT 33.055 384.61 33.255 385.34 ;
      RECT 33.71 384.61 33.91 385.34 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 384.61 34.48 385.34 ;
      RECT 34.775 384.61 34.975 385.34 ;
      RECT 35.27 384.61 35.63 385.34 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 384.61 36.04 385.34 ;
      RECT 36.495 384.61 36.695 385.34 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 384.61 37.265 385.34 ;
      RECT 37.475 384.61 37.675 385.34 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 384.61 38.33 385.34 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 384.61 38.9 385.34 ;
      RECT 39.195 384.61 39.395 385.34 ;
      RECT 39.69 384.61 40.05 385.34 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 384.61 40.46 385.34 ;
      RECT 40.915 384.61 41.115 385.34 ;
      RECT 41.325 384.61 41.685 385.34 ;
      RECT 41.895 384.61 42.095 385.34 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 384.61 42.75 385.34 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 384.61 43.32 385.34 ;
      RECT 43.615 384.61 43.815 385.34 ;
      RECT 44.11 384.61 44.47 385.34 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 384.61 44.88 385.34 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 384.61 45.535 385.34 ;
      RECT 45.745 384.61 46.105 385.34 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 384.61 46.515 385.34 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 384.61 47.17 385.34 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 384.61 47.74 385.34 ;
      RECT 48.035 384.61 48.235 385.34 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 384.61 48.89 385.34 ;
      RECT 49.1 384.61 49.3 385.34 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 384.61 49.955 385.34 ;
      RECT 50.165 384.61 50.525 385.34 ;
      RECT 50.735 384.61 50.935 385.34 ;
      RECT 51.39 384.61 51.59 385.34 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 384.61 52.16 385.34 ;
      RECT 52.455 384.61 52.655 385.34 ;
      RECT 52.95 384.61 53.31 385.34 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 384.61 53.72 385.34 ;
      RECT 54.175 384.61 54.375 385.34 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 384.61 54.945 385.34 ;
      RECT 55.155 384.61 55.355 385.34 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 384.61 56.01 385.34 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 384.61 56.58 385.34 ;
      RECT 56.875 384.61 57.075 385.34 ;
      RECT 57.37 384.61 57.73 385.34 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 384.61 58.14 385.34 ;
      RECT 58.595 384.61 58.795 385.34 ;
      RECT 59.005 384.61 59.365 385.34 ;
      RECT 59.575 384.61 59.775 385.34 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 384.61 60.43 385.34 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 384.61 61 385.34 ;
      RECT 61.295 384.61 61.495 385.34 ;
      RECT 61.79 384.61 62.15 385.34 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 384.61 62.56 385.34 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 384.61 63.215 385.34 ;
      RECT 63.425 384.61 63.785 385.34 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 384.61 64.195 385.34 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 384.61 64.85 385.34 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 384.61 65.42 385.34 ;
      RECT 65.715 384.61 65.915 385.34 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 384.61 66.57 385.34 ;
      RECT 66.78 384.61 66.98 385.34 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 384.61 67.635 385.34 ;
      RECT 67.845 384.61 68.205 385.34 ;
      RECT 68.415 384.61 68.615 385.34 ;
      RECT 69.07 384.61 69.27 385.34 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 384.61 69.84 385.34 ;
      RECT 70.135 384.61 70.335 385.34 ;
      RECT 70.63 384.61 70.99 385.34 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 384.61 71.4 385.34 ;
      RECT 71.855 384.61 72.055 385.34 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 72.265 384.61 72.625 385.34 ;
      RECT 72.835 384.61 73.035 385.34 ;
      RECT 72.91 0.52 73.17 7.78 ;
      RECT 73.42 0.3 73.68 5.235 ;
      RECT 73.49 384.61 73.69 385.34 ;
      RECT 73.93 0.52 74.19 5.57 ;
      RECT 73.9 384.61 74.26 385.34 ;
      RECT 74.555 384.61 74.755 385.34 ;
      RECT 75.05 384.61 75.41 385.34 ;
      RECT 75.305 0.52 75.565 6.28 ;
      RECT 75.62 384.61 75.82 385.34 ;
      RECT 76.275 384.61 76.475 385.34 ;
      RECT 76.685 384.61 77.045 385.34 ;
      RECT 77.255 384.61 77.455 385.34 ;
      RECT 76.99 0.18 77.76 0.88 ;
      RECT 77.91 384.61 78.11 385.34 ;
      RECT 78.01 0.3 78.27 8.7 ;
      RECT 78.32 384.61 78.68 385.34 ;
      RECT 78.975 384.61 79.175 385.34 ;
      RECT 79.47 384.61 79.83 385.34 ;
      RECT 80.56 0.155 81.33 0.445 ;
      RECT 80.56 0.155 80.82 8.665 ;
      RECT 81.07 0.155 81.33 8.665 ;
      RECT 80.04 384.61 80.24 385.34 ;
      RECT 80.05 0.52 80.31 9.955 ;
      RECT 80.695 384.61 80.895 385.34 ;
      RECT 81.105 384.61 81.465 385.34 ;
      RECT 81.58 0.52 81.84 11.315 ;
      RECT 81.675 384.61 81.875 385.34 ;
      RECT 82.09 0.52 82.35 13.45 ;
      RECT 82.33 384.61 82.53 385.34 ;
      RECT 82.6 0.52 82.86 14.115 ;
      RECT 82.74 384.61 83.1 385.34 ;
      RECT 83.395 384.61 83.595 385.34 ;
      RECT 84.795 0.155 85.565 0.445 ;
      RECT 84.795 0.155 85.055 13.21 ;
      RECT 85.305 0.155 85.565 13.21 ;
      RECT 83.89 384.61 84.25 385.34 ;
      RECT 84.46 384.61 84.66 385.34 ;
      RECT 85.815 0.18 86.585 0.88 ;
      RECT 85.815 0.18 86.075 12.9 ;
      RECT 86.325 0.18 86.585 12.9 ;
      RECT 85.115 384.61 85.315 385.34 ;
      RECT 85.525 384.61 85.885 385.34 ;
      RECT 86.095 384.61 86.295 385.34 ;
      RECT 86.75 384.61 86.95 385.34 ;
      RECT 87.035 0.52 87.295 2.82 ;
      RECT 87.16 384.61 87.52 385.34 ;
      RECT 87.815 384.61 88.015 385.34 ;
      RECT 88.31 384.61 88.67 385.34 ;
      RECT 88.565 0.52 88.825 2.82 ;
      RECT 88.88 384.61 89.08 385.34 ;
      RECT 89.535 384.61 89.735 385.34 ;
      RECT 89.74 0.52 90 4.315 ;
      RECT 89.945 384.61 90.305 385.34 ;
      RECT 90.515 384.61 90.715 385.34 ;
      RECT 90.59 0.52 90.85 7.78 ;
      RECT 91.1 0.3 91.36 5.235 ;
      RECT 91.17 384.61 91.37 385.34 ;
      RECT 91.61 0.52 91.87 5.57 ;
      RECT 91.58 384.61 91.94 385.34 ;
      RECT 92.235 384.61 92.435 385.34 ;
      RECT 92.73 384.61 93.09 385.34 ;
      RECT 92.985 0.52 93.245 6.28 ;
      RECT 93.3 384.61 93.5 385.34 ;
      RECT 93.955 384.61 94.155 385.34 ;
      RECT 94.365 384.61 94.725 385.34 ;
      RECT 94.935 384.61 95.135 385.34 ;
      RECT 94.67 0.18 95.44 0.88 ;
      RECT 95.59 384.61 95.79 385.34 ;
      RECT 95.69 0.3 95.95 8.7 ;
      RECT 96 384.61 96.36 385.34 ;
      RECT 96.655 384.61 96.855 385.34 ;
      RECT 97.15 384.61 97.51 385.34 ;
      RECT 98.24 0.155 99.01 0.445 ;
      RECT 98.24 0.155 98.5 8.665 ;
      RECT 98.75 0.155 99.01 8.665 ;
      RECT 97.72 384.61 97.92 385.34 ;
      RECT 97.73 0.52 97.99 9.955 ;
      RECT 98.375 384.61 98.575 385.34 ;
      RECT 98.785 384.61 99.145 385.34 ;
      RECT 99.26 0.52 99.52 11.315 ;
      RECT 99.355 384.61 99.555 385.34 ;
      RECT 99.77 0.52 100.03 13.45 ;
      RECT 100.01 384.61 100.21 385.34 ;
      RECT 100.28 0.52 100.54 14.115 ;
      RECT 100.42 384.61 100.78 385.34 ;
      RECT 101.075 384.61 101.275 385.34 ;
      RECT 102.475 0.155 103.245 0.445 ;
      RECT 102.475 0.155 102.735 13.21 ;
      RECT 102.985 0.155 103.245 13.21 ;
      RECT 101.57 384.61 101.93 385.34 ;
      RECT 102.14 384.61 102.34 385.34 ;
      RECT 103.495 0.18 104.265 0.88 ;
      RECT 103.495 0.18 103.755 12.9 ;
      RECT 104.005 0.18 104.265 12.9 ;
      RECT 102.795 384.61 102.995 385.34 ;
      RECT 103.205 384.61 103.565 385.34 ;
      RECT 103.775 384.61 103.975 385.34 ;
      RECT 104.43 384.61 104.63 385.34 ;
      RECT 104.715 0.52 104.975 2.82 ;
      RECT 104.84 384.61 105.2 385.34 ;
      RECT 105.495 384.61 105.695 385.34 ;
      RECT 105.99 384.61 106.35 385.34 ;
      RECT 106.245 0.52 106.505 2.82 ;
      RECT 106.56 384.61 106.76 385.34 ;
      RECT 107.215 384.61 107.415 385.34 ;
      RECT 107.42 0.52 107.68 4.315 ;
      RECT 107.625 384.61 107.985 385.34 ;
      RECT 108.195 384.61 108.395 385.34 ;
      RECT 108.27 0.52 108.53 7.78 ;
      RECT 108.78 0.3 109.04 5.235 ;
      RECT 108.85 384.61 109.05 385.34 ;
      RECT 109.29 0.52 109.55 5.57 ;
      RECT 109.26 384.61 109.62 385.34 ;
      RECT 109.915 384.61 110.115 385.34 ;
      RECT 110.41 384.61 110.77 385.34 ;
      RECT 110.665 0.52 110.925 6.28 ;
      RECT 110.98 384.61 111.18 385.34 ;
      RECT 111.635 384.61 111.835 385.34 ;
      RECT 112.045 384.61 112.405 385.34 ;
      RECT 112.615 384.61 112.815 385.34 ;
      RECT 112.35 0.18 113.12 0.88 ;
      RECT 113.27 384.61 113.47 385.34 ;
      RECT 113.37 0.3 113.63 8.7 ;
      RECT 113.68 384.61 114.04 385.34 ;
      RECT 114.335 384.61 114.535 385.34 ;
      RECT 114.83 384.61 115.19 385.34 ;
      RECT 115.92 0.155 116.69 0.445 ;
      RECT 115.92 0.155 116.18 8.665 ;
      RECT 116.43 0.155 116.69 8.665 ;
      RECT 115.4 384.61 115.6 385.34 ;
      RECT 115.41 0.52 115.67 9.955 ;
      RECT 116.055 384.61 116.255 385.34 ;
      RECT 116.465 384.61 116.825 385.34 ;
      RECT 116.94 0.52 117.2 11.315 ;
      RECT 117.035 384.61 117.235 385.34 ;
      RECT 117.45 0.52 117.71 13.45 ;
      RECT 117.69 384.61 117.89 385.34 ;
      RECT 117.96 0.52 118.22 14.115 ;
      RECT 118.1 384.61 118.46 385.34 ;
      RECT 118.755 384.61 118.955 385.34 ;
      RECT 120.155 0.155 120.925 0.445 ;
      RECT 120.155 0.155 120.415 13.21 ;
      RECT 120.665 0.155 120.925 13.21 ;
      RECT 119.25 384.61 119.61 385.34 ;
      RECT 119.82 384.61 120.02 385.34 ;
      RECT 121.175 0.18 121.945 0.88 ;
      RECT 121.175 0.18 121.435 12.9 ;
      RECT 121.685 0.18 121.945 12.9 ;
      RECT 120.475 384.61 120.675 385.34 ;
      RECT 120.885 384.61 121.245 385.34 ;
      RECT 121.455 384.61 121.655 385.34 ;
      RECT 122.11 384.61 122.31 385.34 ;
      RECT 122.395 0.52 122.655 2.82 ;
      RECT 122.52 384.61 122.88 385.34 ;
      RECT 123.175 384.61 123.375 385.34 ;
      RECT 123.67 384.61 124.03 385.34 ;
      RECT 123.925 0.52 124.185 2.82 ;
      RECT 124.24 384.61 124.44 385.34 ;
      RECT 124.895 384.61 125.095 385.34 ;
      RECT 125.1 0.52 125.36 4.315 ;
      RECT 125.305 384.61 125.665 385.34 ;
      RECT 125.875 384.61 126.075 385.34 ;
      RECT 125.95 0.52 126.21 7.78 ;
      RECT 126.46 0.3 126.72 5.235 ;
      RECT 126.53 384.61 126.73 385.34 ;
      RECT 126.97 0.52 127.23 5.57 ;
      RECT 126.94 384.61 127.3 385.34 ;
      RECT 127.595 384.61 127.795 385.34 ;
      RECT 128.09 384.61 128.45 385.34 ;
      RECT 128.345 0.52 128.605 6.28 ;
      RECT 128.66 384.61 128.86 385.34 ;
      RECT 129.315 384.61 129.515 385.34 ;
      RECT 129.725 384.61 130.085 385.34 ;
      RECT 130.295 384.61 130.495 385.34 ;
      RECT 130.03 0.18 130.8 0.88 ;
      RECT 130.95 384.61 131.15 385.34 ;
      RECT 131.05 0.3 131.31 8.7 ;
      RECT 131.36 384.61 131.72 385.34 ;
      RECT 132.015 384.61 132.215 385.34 ;
      RECT 132.51 384.61 132.87 385.34 ;
      RECT 133.6 0.155 134.37 0.445 ;
      RECT 133.6 0.155 133.86 8.665 ;
      RECT 134.11 0.155 134.37 8.665 ;
      RECT 133.08 384.61 133.28 385.34 ;
      RECT 133.09 0.52 133.35 9.955 ;
      RECT 133.735 384.61 133.935 385.34 ;
      RECT 134.145 384.61 134.505 385.34 ;
      RECT 134.62 0.52 134.88 11.315 ;
      RECT 134.715 384.61 134.915 385.34 ;
      RECT 135.13 0.52 135.39 13.45 ;
      RECT 135.37 384.61 135.57 385.34 ;
      RECT 135.64 0.52 135.9 14.115 ;
      RECT 135.78 384.61 136.14 385.34 ;
      RECT 136.435 384.61 136.635 385.34 ;
      RECT 137.835 0.155 138.605 0.445 ;
      RECT 137.835 0.155 138.095 13.21 ;
      RECT 138.345 0.155 138.605 13.21 ;
      RECT 136.93 384.61 137.29 385.34 ;
      RECT 137.5 384.61 137.7 385.34 ;
      RECT 138.855 0.18 139.625 0.88 ;
      RECT 138.855 0.18 139.115 12.9 ;
      RECT 139.365 0.18 139.625 12.9 ;
      RECT 138.155 384.61 138.355 385.34 ;
      RECT 138.565 384.61 138.925 385.34 ;
      RECT 139.135 384.61 139.335 385.34 ;
      RECT 139.79 384.61 139.99 385.34 ;
      RECT 140.075 0.52 140.335 2.82 ;
      RECT 140.2 384.61 140.56 385.34 ;
      RECT 140.855 384.61 141.055 385.34 ;
      RECT 141.35 384.61 141.71 385.34 ;
      RECT 141.605 0.52 141.865 2.82 ;
      RECT 141.92 384.61 142.12 385.34 ;
      RECT 142.575 384.61 142.775 385.34 ;
      RECT 142.78 0.52 143.04 4.315 ;
      RECT 142.985 384.61 143.345 385.34 ;
      RECT 143.555 384.61 143.755 385.34 ;
      RECT 143.63 0.52 143.89 7.78 ;
      RECT 144.14 0.3 144.4 5.235 ;
      RECT 144.21 384.61 144.41 385.34 ;
      RECT 144.65 0.52 144.91 5.57 ;
      RECT 144.62 384.61 144.98 385.34 ;
      RECT 145.275 384.61 145.475 385.34 ;
      RECT 145.77 384.61 146.13 385.34 ;
      RECT 146.025 0.52 146.285 6.28 ;
      RECT 146.34 384.61 146.54 385.34 ;
      RECT 146.995 384.61 147.195 385.34 ;
      RECT 147.405 384.61 147.765 385.34 ;
      RECT 147.975 384.61 148.175 385.34 ;
      RECT 147.71 0.18 148.48 0.88 ;
      RECT 148.63 384.61 148.83 385.34 ;
      RECT 148.73 0.3 148.99 8.7 ;
      RECT 149.04 384.61 149.4 385.34 ;
      RECT 149.695 384.61 149.895 385.34 ;
      RECT 150.19 384.61 150.55 385.34 ;
      RECT 151.28 0.155 152.05 0.445 ;
      RECT 151.28 0.155 151.54 8.665 ;
      RECT 151.79 0.155 152.05 8.665 ;
      RECT 150.76 384.61 150.96 385.34 ;
      RECT 150.77 0.52 151.03 9.955 ;
      RECT 151.415 384.61 151.615 385.34 ;
      RECT 151.825 384.61 152.185 385.34 ;
      RECT 152.3 0.52 152.56 11.315 ;
      RECT 152.395 384.61 152.595 385.34 ;
      RECT 152.81 0.52 153.07 13.45 ;
      RECT 153.05 384.61 153.25 385.34 ;
      RECT 153.32 0.52 153.58 14.115 ;
      RECT 153.46 384.61 153.82 385.34 ;
      RECT 154.115 384.61 154.315 385.34 ;
      RECT 155.515 0.155 156.285 0.445 ;
      RECT 155.515 0.155 155.775 13.21 ;
      RECT 156.025 0.155 156.285 13.21 ;
      RECT 154.61 384.61 154.97 385.34 ;
      RECT 155.18 384.61 155.38 385.34 ;
      RECT 156.535 0.18 157.305 0.88 ;
      RECT 156.535 0.18 156.795 12.9 ;
      RECT 157.045 0.18 157.305 12.9 ;
      RECT 155.835 384.61 156.035 385.34 ;
      RECT 156.245 384.61 156.605 385.34 ;
      RECT 156.815 384.61 157.015 385.34 ;
      RECT 157.47 384.61 157.67 385.34 ;
      RECT 157.755 0.52 158.015 2.82 ;
      RECT 157.88 384.61 158.24 385.34 ;
      RECT 158.535 384.61 158.735 385.34 ;
      RECT 159.03 384.61 159.39 385.34 ;
      RECT 159.285 0.52 159.545 2.82 ;
      RECT 159.6 384.61 159.8 385.34 ;
      RECT 160.255 384.61 160.455 385.34 ;
      RECT 160.46 0.52 160.72 4.315 ;
      RECT 160.665 384.61 161.025 385.34 ;
      RECT 161.235 384.61 161.435 385.34 ;
      RECT 161.31 0.52 161.57 7.78 ;
      RECT 161.82 0.3 162.08 5.235 ;
      RECT 161.89 384.61 162.09 385.34 ;
      RECT 162.33 0.52 162.59 5.57 ;
      RECT 162.3 384.61 162.66 385.34 ;
      RECT 162.955 384.61 163.155 385.34 ;
      RECT 163.45 384.61 163.81 385.34 ;
      RECT 163.705 0.52 163.965 6.28 ;
      RECT 164.02 384.61 164.22 385.34 ;
      RECT 164.675 384.61 164.875 385.34 ;
      RECT 165.085 384.61 165.445 385.34 ;
      RECT 165.655 384.61 165.855 385.34 ;
      RECT 165.39 0.18 166.16 0.88 ;
      RECT 166.31 384.61 166.51 385.34 ;
      RECT 166.41 0.3 166.67 8.7 ;
      RECT 166.72 384.61 167.08 385.34 ;
      RECT 167.375 384.61 167.575 385.34 ;
      RECT 167.87 384.61 168.23 385.34 ;
      RECT 168.96 0.155 169.73 0.445 ;
      RECT 168.96 0.155 169.22 8.665 ;
      RECT 169.47 0.155 169.73 8.665 ;
      RECT 168.44 384.61 168.64 385.34 ;
      RECT 168.45 0.52 168.71 9.955 ;
      RECT 169.095 384.61 169.295 385.34 ;
      RECT 169.505 384.61 169.865 385.34 ;
      RECT 169.98 0.52 170.24 11.315 ;
      RECT 170.075 384.61 170.275 385.34 ;
      RECT 170.49 0.52 170.75 13.45 ;
      RECT 170.73 384.61 170.93 385.34 ;
      RECT 171 0.52 171.26 14.115 ;
      RECT 171.14 384.61 171.5 385.34 ;
      RECT 171.795 384.61 171.995 385.34 ;
      RECT 173.195 0.155 173.965 0.445 ;
      RECT 173.195 0.155 173.455 13.21 ;
      RECT 173.705 0.155 173.965 13.21 ;
      RECT 172.29 384.61 172.65 385.34 ;
      RECT 172.86 384.61 173.06 385.34 ;
      RECT 174.215 0.18 174.985 0.88 ;
      RECT 174.215 0.18 174.475 12.9 ;
      RECT 174.725 0.18 174.985 12.9 ;
      RECT 173.515 384.61 173.715 385.34 ;
      RECT 173.925 384.61 174.285 385.34 ;
      RECT 174.495 384.61 174.695 385.34 ;
      RECT 175.15 384.61 175.35 385.34 ;
      RECT 175.435 0.52 175.695 2.82 ;
      RECT 175.56 384.61 175.92 385.34 ;
      RECT 176.215 384.61 176.415 385.34 ;
      RECT 176.71 384.61 177.07 385.34 ;
      RECT 176.965 0.52 177.225 2.82 ;
      RECT 177.28 384.61 177.48 385.34 ;
      RECT 177.935 384.61 178.135 385.34 ;
      RECT 178.14 0.52 178.4 4.315 ;
      RECT 178.345 384.61 178.705 385.34 ;
      RECT 178.915 384.61 179.115 385.34 ;
      RECT 178.99 0.52 179.25 7.78 ;
      RECT 179.5 0.3 179.76 5.235 ;
      RECT 179.57 384.61 179.77 385.34 ;
      RECT 180.01 0.52 180.27 5.57 ;
      RECT 179.98 384.61 180.34 385.34 ;
      RECT 180.635 384.61 180.835 385.34 ;
      RECT 181.13 384.61 181.49 385.34 ;
      RECT 181.385 0.52 181.645 6.28 ;
      RECT 181.7 384.61 181.9 385.34 ;
      RECT 182.355 384.61 182.555 385.34 ;
      RECT 182.765 384.61 183.125 385.34 ;
      RECT 183.335 384.61 183.535 385.34 ;
      RECT 183.07 0.18 183.84 0.88 ;
      RECT 183.99 384.61 184.19 385.34 ;
      RECT 184.09 0.3 184.35 8.7 ;
      RECT 184.4 384.61 184.76 385.34 ;
      RECT 185.055 384.61 185.255 385.34 ;
      RECT 185.55 384.61 185.91 385.34 ;
      RECT 186.64 0.155 187.41 0.445 ;
      RECT 186.64 0.155 186.9 8.665 ;
      RECT 187.15 0.155 187.41 8.665 ;
      RECT 186.12 384.61 186.32 385.34 ;
      RECT 186.13 0.52 186.39 9.955 ;
      RECT 186.775 384.61 186.975 385.34 ;
      RECT 187.185 384.61 187.545 385.34 ;
      RECT 187.66 0.52 187.92 11.315 ;
      RECT 187.755 384.61 187.955 385.34 ;
      RECT 188.17 0.52 188.43 13.45 ;
      RECT 188.41 384.61 188.61 385.34 ;
      RECT 188.68 0.52 188.94 14.115 ;
      RECT 188.82 384.61 189.18 385.34 ;
      RECT 189.475 384.61 189.675 385.34 ;
      RECT 190.875 0.155 191.645 0.445 ;
      RECT 190.875 0.155 191.135 13.21 ;
      RECT 191.385 0.155 191.645 13.21 ;
      RECT 189.97 384.61 190.33 385.34 ;
      RECT 190.54 384.61 190.74 385.34 ;
      RECT 191.895 0.18 192.665 0.88 ;
      RECT 191.895 0.18 192.155 12.9 ;
      RECT 192.405 0.18 192.665 12.9 ;
      RECT 191.195 384.61 191.395 385.34 ;
      RECT 191.605 384.61 191.965 385.34 ;
      RECT 192.175 384.61 192.375 385.34 ;
      RECT 192.83 384.61 193.03 385.34 ;
      RECT 193.115 0.52 193.375 2.82 ;
      RECT 193.24 384.61 193.6 385.34 ;
      RECT 193.895 384.61 194.095 385.34 ;
      RECT 194.39 384.61 194.75 385.34 ;
      RECT 194.645 0.52 194.905 2.82 ;
      RECT 194.96 384.61 195.16 385.34 ;
      RECT 195.615 384.61 195.815 385.34 ;
      RECT 195.82 0.52 196.08 4.315 ;
      RECT 196.025 384.61 196.385 385.34 ;
      RECT 196.595 384.61 196.795 385.34 ;
      RECT 196.67 0.52 196.93 7.78 ;
      RECT 197.18 0.3 197.44 5.235 ;
      RECT 197.25 384.61 197.45 385.34 ;
      RECT 197.69 0.52 197.95 5.57 ;
      RECT 197.66 384.61 198.02 385.34 ;
      RECT 198.315 384.61 198.515 385.34 ;
      RECT 198.81 384.61 199.17 385.34 ;
      RECT 199.065 0.52 199.325 6.28 ;
      RECT 199.38 384.61 199.58 385.34 ;
      RECT 200.035 384.61 200.235 385.34 ;
      RECT 200.445 384.61 200.805 385.34 ;
      RECT 201.015 384.61 201.215 385.34 ;
      RECT 200.75 0.18 201.52 0.88 ;
      RECT 201.67 384.61 201.87 385.34 ;
      RECT 201.77 0.3 202.03 8.7 ;
      RECT 202.08 384.61 202.44 385.34 ;
      RECT 202.735 384.61 202.935 385.34 ;
      RECT 203.23 384.61 203.59 385.34 ;
      RECT 204.32 0.155 205.09 0.445 ;
      RECT 204.32 0.155 204.58 8.665 ;
      RECT 204.83 0.155 205.09 8.665 ;
      RECT 203.8 384.61 204 385.34 ;
      RECT 203.81 0.52 204.07 9.955 ;
      RECT 204.455 384.61 204.655 385.34 ;
      RECT 204.865 384.61 205.225 385.34 ;
      RECT 205.34 0.52 205.6 11.315 ;
      RECT 205.435 384.61 205.635 385.34 ;
      RECT 205.85 0.52 206.11 13.45 ;
      RECT 206.09 384.61 206.29 385.34 ;
      RECT 206.36 0.52 206.62 14.115 ;
      RECT 206.5 384.61 206.86 385.34 ;
      RECT 207.155 384.61 207.355 385.34 ;
      RECT 208.555 0.155 209.325 0.445 ;
      RECT 208.555 0.155 208.815 13.21 ;
      RECT 209.065 0.155 209.325 13.21 ;
      RECT 207.65 384.61 208.01 385.34 ;
      RECT 208.22 384.61 208.42 385.34 ;
      RECT 209.575 0.18 210.345 0.88 ;
      RECT 209.575 0.18 209.835 12.9 ;
      RECT 210.085 0.18 210.345 12.9 ;
      RECT 208.875 384.61 209.075 385.34 ;
      RECT 209.285 384.61 209.645 385.34 ;
      RECT 209.855 384.61 210.055 385.34 ;
      RECT 210.51 384.61 210.71 385.34 ;
      RECT 210.795 0.52 211.055 2.82 ;
      RECT 210.92 384.61 211.28 385.34 ;
      RECT 211.575 384.61 211.775 385.34 ;
      RECT 212.07 384.61 212.43 385.34 ;
      RECT 212.325 0.52 212.585 2.82 ;
      RECT 212.64 384.61 212.84 385.34 ;
      RECT 213.295 384.61 213.495 385.34 ;
      RECT 213.5 0.52 213.76 4.315 ;
      RECT 213.705 384.61 214.065 385.34 ;
      RECT 214.275 384.61 214.475 385.34 ;
      RECT 214.35 0.52 214.61 7.78 ;
      RECT 214.86 0.3 215.12 5.235 ;
      RECT 214.93 384.61 215.13 385.34 ;
      RECT 215.37 0.52 215.63 5.57 ;
      RECT 215.34 384.61 215.7 385.34 ;
      RECT 215.995 384.61 216.195 385.34 ;
      RECT 216.49 384.61 216.85 385.34 ;
      RECT 216.745 0.52 217.005 6.28 ;
      RECT 217.06 384.61 217.26 385.34 ;
      RECT 217.715 384.61 217.915 385.34 ;
      RECT 218.125 384.61 218.485 385.34 ;
      RECT 218.695 384.61 218.895 385.34 ;
      RECT 218.43 0.18 219.2 0.88 ;
      RECT 219.35 384.61 219.55 385.34 ;
      RECT 219.45 0.3 219.71 8.7 ;
      RECT 219.76 384.61 220.12 385.34 ;
      RECT 220.415 384.61 220.615 385.34 ;
      RECT 220.91 384.61 221.27 385.34 ;
      RECT 222 0.155 222.77 0.445 ;
      RECT 222 0.155 222.26 8.665 ;
      RECT 222.51 0.155 222.77 8.665 ;
      RECT 221.48 384.61 221.68 385.34 ;
      RECT 221.49 0.52 221.75 9.955 ;
      RECT 222.135 384.61 222.335 385.34 ;
      RECT 222.545 384.61 222.905 385.34 ;
      RECT 223.02 0.52 223.28 11.315 ;
      RECT 223.115 384.61 223.315 385.34 ;
      RECT 223.53 0.52 223.79 13.45 ;
      RECT 223.77 384.61 223.97 385.34 ;
      RECT 224.04 0.52 224.3 14.115 ;
      RECT 224.18 384.61 224.54 385.34 ;
      RECT 224.835 384.61 225.035 385.34 ;
      RECT 226.235 0.155 227.005 0.445 ;
      RECT 226.235 0.155 226.495 13.21 ;
      RECT 226.745 0.155 227.005 13.21 ;
      RECT 225.33 384.61 225.69 385.34 ;
      RECT 225.9 384.61 226.1 385.34 ;
      RECT 227.255 0.18 228.025 0.88 ;
      RECT 227.255 0.18 227.515 12.9 ;
      RECT 227.765 0.18 228.025 12.9 ;
      RECT 226.555 384.61 226.755 385.34 ;
      RECT 226.965 384.61 227.325 385.34 ;
      RECT 227.535 384.61 227.735 385.34 ;
      RECT 228.19 384.61 228.39 385.34 ;
      RECT 228.475 0.52 228.735 2.82 ;
      RECT 228.6 384.61 228.96 385.34 ;
      RECT 229.255 384.61 229.455 385.34 ;
      RECT 229.75 384.61 230.11 385.34 ;
      RECT 230.005 0.52 230.265 2.82 ;
      RECT 230.32 384.61 230.52 385.34 ;
      RECT 230.975 384.61 231.175 385.34 ;
      RECT 231.18 0.52 231.44 4.315 ;
      RECT 231.385 384.61 231.745 385.34 ;
      RECT 231.955 384.61 232.155 385.34 ;
      RECT 232.03 0.52 232.29 7.78 ;
      RECT 232.54 0.3 232.8 5.235 ;
      RECT 232.61 384.61 232.81 385.34 ;
      RECT 233.05 0.52 233.31 5.57 ;
      RECT 233.02 384.61 233.38 385.34 ;
      RECT 233.675 384.61 233.875 385.34 ;
      RECT 234.17 384.61 234.53 385.34 ;
      RECT 234.425 0.52 234.685 6.28 ;
      RECT 234.74 384.61 234.94 385.34 ;
      RECT 235.395 384.61 235.595 385.34 ;
      RECT 235.805 384.61 236.165 385.34 ;
      RECT 236.375 384.61 236.575 385.34 ;
      RECT 236.11 0.18 236.88 0.88 ;
      RECT 237.03 384.61 237.23 385.34 ;
      RECT 237.13 0.3 237.39 8.7 ;
      RECT 237.44 384.61 237.8 385.34 ;
      RECT 238.095 384.61 238.295 385.34 ;
      RECT 238.59 384.61 238.95 385.34 ;
      RECT 239.68 0.155 240.45 0.445 ;
      RECT 239.68 0.155 239.94 8.665 ;
      RECT 240.19 0.155 240.45 8.665 ;
      RECT 239.16 384.61 239.36 385.34 ;
      RECT 239.17 0.52 239.43 9.955 ;
      RECT 239.815 384.61 240.015 385.34 ;
      RECT 240.225 384.61 240.585 385.34 ;
      RECT 240.7 0.52 240.96 11.315 ;
      RECT 240.795 384.61 240.995 385.34 ;
      RECT 241.21 0.52 241.47 13.45 ;
      RECT 241.45 384.61 241.65 385.34 ;
      RECT 241.72 0.52 241.98 14.115 ;
      RECT 241.86 384.61 242.22 385.34 ;
      RECT 242.515 384.61 242.715 385.34 ;
      RECT 243.915 0.155 244.685 0.445 ;
      RECT 243.915 0.155 244.175 13.21 ;
      RECT 244.425 0.155 244.685 13.21 ;
      RECT 243.01 384.61 243.37 385.34 ;
      RECT 243.58 384.61 243.78 385.34 ;
      RECT 244.935 0.18 245.705 0.88 ;
      RECT 244.935 0.18 245.195 12.9 ;
      RECT 245.445 0.18 245.705 12.9 ;
      RECT 244.235 384.61 244.435 385.34 ;
      RECT 244.645 384.61 245.005 385.34 ;
      RECT 245.215 384.61 245.415 385.34 ;
      RECT 245.87 384.61 246.07 385.34 ;
      RECT 246.155 0.52 246.415 2.82 ;
      RECT 246.28 384.61 246.64 385.34 ;
      RECT 246.935 384.61 247.135 385.34 ;
      RECT 247.43 384.61 247.79 385.34 ;
      RECT 247.685 0.52 247.945 2.82 ;
      RECT 248 384.61 248.2 385.34 ;
      RECT 248.655 384.61 248.855 385.34 ;
      RECT 248.86 0.52 249.12 4.315 ;
      RECT 249.065 384.61 249.425 385.34 ;
      RECT 249.635 384.61 249.835 385.34 ;
      RECT 249.71 0.52 249.97 7.78 ;
      RECT 250.22 0.3 250.48 5.235 ;
      RECT 250.29 384.61 250.49 385.34 ;
      RECT 250.73 0.52 250.99 5.57 ;
      RECT 250.7 384.61 251.06 385.34 ;
      RECT 251.355 384.61 251.555 385.34 ;
      RECT 251.85 384.61 252.21 385.34 ;
      RECT 252.105 0.52 252.365 6.28 ;
      RECT 252.42 384.61 252.62 385.34 ;
      RECT 253.075 384.61 253.275 385.34 ;
      RECT 253.485 384.61 253.845 385.34 ;
      RECT 254.055 384.61 254.255 385.34 ;
      RECT 253.79 0.18 254.56 0.88 ;
      RECT 254.71 384.61 254.91 385.34 ;
      RECT 254.81 0.3 255.07 8.7 ;
      RECT 255.12 384.61 255.48 385.34 ;
      RECT 255.775 384.61 255.975 385.34 ;
      RECT 256.27 384.61 256.63 385.34 ;
      RECT 257.36 0.155 258.13 0.445 ;
      RECT 257.36 0.155 257.62 8.665 ;
      RECT 257.87 0.155 258.13 8.665 ;
      RECT 256.84 384.61 257.04 385.34 ;
      RECT 256.85 0.52 257.11 9.955 ;
      RECT 257.495 384.61 257.695 385.34 ;
      RECT 257.905 384.61 258.265 385.34 ;
      RECT 258.38 0.52 258.64 11.315 ;
      RECT 258.475 384.61 258.675 385.34 ;
      RECT 258.89 0.52 259.15 13.45 ;
      RECT 259.13 384.61 259.33 385.34 ;
      RECT 259.4 0.52 259.66 14.115 ;
      RECT 259.54 384.61 259.9 385.34 ;
      RECT 260.195 384.61 260.395 385.34 ;
      RECT 261.595 0.155 262.365 0.445 ;
      RECT 261.595 0.155 261.855 13.21 ;
      RECT 262.105 0.155 262.365 13.21 ;
      RECT 260.69 384.61 261.05 385.34 ;
      RECT 261.26 384.61 261.46 385.34 ;
      RECT 262.615 0.18 263.385 0.88 ;
      RECT 262.615 0.18 262.875 12.9 ;
      RECT 263.125 0.18 263.385 12.9 ;
      RECT 261.915 384.61 262.115 385.34 ;
      RECT 262.325 384.61 262.685 385.34 ;
      RECT 262.895 384.61 263.095 385.34 ;
      RECT 263.55 384.61 263.75 385.34 ;
      RECT 263.835 0.52 264.095 2.82 ;
      RECT 263.96 384.61 264.32 385.34 ;
      RECT 264.615 384.61 264.815 385.34 ;
      RECT 265.11 384.61 265.47 385.34 ;
      RECT 265.365 0.52 265.625 2.82 ;
      RECT 265.68 384.61 265.88 385.34 ;
      RECT 266.335 384.61 266.535 385.34 ;
      RECT 266.54 0.52 266.8 4.315 ;
      RECT 266.745 384.61 267.105 385.34 ;
      RECT 267.315 384.61 267.515 385.34 ;
      RECT 267.39 0.52 267.65 7.78 ;
      RECT 267.9 0.3 268.16 5.235 ;
      RECT 267.97 384.61 268.17 385.34 ;
      RECT 268.41 0.52 268.67 5.57 ;
      RECT 268.38 384.61 268.74 385.34 ;
      RECT 269.035 384.61 269.235 385.34 ;
      RECT 269.53 384.61 269.89 385.34 ;
      RECT 269.785 0.52 270.045 6.28 ;
      RECT 270.1 384.61 270.3 385.34 ;
      RECT 270.755 384.61 270.955 385.34 ;
      RECT 271.165 384.61 271.525 385.34 ;
      RECT 271.735 384.61 271.935 385.34 ;
      RECT 271.47 0.18 272.24 0.88 ;
      RECT 272.39 384.61 272.59 385.34 ;
      RECT 272.49 0.3 272.75 8.7 ;
      RECT 272.8 384.61 273.16 385.34 ;
      RECT 273.455 384.61 273.655 385.34 ;
      RECT 273.95 384.61 274.31 385.34 ;
      RECT 275.04 0.155 275.81 0.445 ;
      RECT 275.04 0.155 275.3 8.665 ;
      RECT 275.55 0.155 275.81 8.665 ;
      RECT 274.52 384.61 274.72 385.34 ;
      RECT 274.53 0.52 274.79 9.955 ;
      RECT 275.175 384.61 275.375 385.34 ;
      RECT 275.585 384.61 275.945 385.34 ;
      RECT 276.06 0.52 276.32 11.315 ;
      RECT 276.155 384.61 276.355 385.34 ;
      RECT 276.57 0.52 276.83 13.45 ;
      RECT 276.81 384.61 277.01 385.34 ;
      RECT 277.08 0.52 277.34 14.115 ;
      RECT 277.22 384.61 277.58 385.34 ;
      RECT 277.875 384.61 278.075 385.34 ;
      RECT 279.275 0.155 280.045 0.445 ;
      RECT 279.275 0.155 279.535 13.21 ;
      RECT 279.785 0.155 280.045 13.21 ;
      RECT 278.37 384.61 278.73 385.34 ;
      RECT 278.94 384.61 279.14 385.34 ;
      RECT 280.295 0.18 281.065 0.88 ;
      RECT 280.295 0.18 280.555 12.9 ;
      RECT 280.805 0.18 281.065 12.9 ;
      RECT 279.595 384.61 279.795 385.34 ;
      RECT 280.005 384.61 280.365 385.34 ;
      RECT 280.575 384.61 280.775 385.34 ;
      RECT 281.23 384.61 281.43 385.34 ;
      RECT 281.515 0.52 281.775 2.82 ;
      RECT 281.64 384.61 282 385.34 ;
      RECT 282.295 384.61 282.495 385.34 ;
      RECT 282.79 384.61 283.15 385.34 ;
      RECT 283.045 0.52 283.305 2.82 ;
      RECT 283.36 384.61 283.56 385.34 ;
      RECT 284.015 384.61 284.215 385.34 ;
      RECT 285.24 0.17 286.01 0.43 ;
      RECT 285.24 0.17 285.5 8.7 ;
      RECT 285.75 0.17 286.01 8.7 ;
      RECT 284.22 0.52 284.48 4.315 ;
      RECT 286.26 0.18 287.03 0.88 ;
      RECT 286.26 0.18 286.52 8.7 ;
      RECT 286.77 0.18 287.03 8.7 ;
      RECT 287.28 0.17 288.05 0.43 ;
      RECT 287.28 0.17 287.54 8.7 ;
      RECT 287.79 0.17 288.05 8.7 ;
      RECT 288.3 0.18 289.07 0.88 ;
      RECT 288.3 0.18 288.56 8.7 ;
      RECT 288.81 0.18 289.07 8.7 ;
      RECT 289.32 0.17 290.09 0.43 ;
      RECT 289.32 0.17 289.58 8.7 ;
      RECT 289.83 0.17 290.09 8.7 ;
      RECT 290.34 0.18 291.11 0.88 ;
      RECT 290.34 0.18 290.6 8.7 ;
      RECT 290.85 0.18 291.11 8.7 ;
      RECT 291.36 0.17 292.13 0.43 ;
      RECT 291.36 0.17 291.62 8.7 ;
      RECT 291.87 0.17 292.13 8.7 ;
      RECT 292.38 0.18 293.15 0.88 ;
      RECT 292.38 0.18 292.64 8.7 ;
      RECT 292.89 0.18 293.15 8.7 ;
      RECT 293.4 0.17 294.17 0.43 ;
      RECT 293.4 0.17 293.66 8.7 ;
      RECT 293.91 0.17 294.17 8.7 ;
      RECT 294.42 0.18 295.19 0.88 ;
      RECT 294.42 0.18 294.68 8.7 ;
      RECT 294.93 0.18 295.19 8.7 ;
      RECT 295.44 0.17 296.21 0.43 ;
      RECT 295.44 0.17 295.7 8.7 ;
      RECT 295.95 0.17 296.21 8.7 ;
      RECT 296.46 0.18 297.23 0.88 ;
      RECT 296.46 0.18 296.72 8.7 ;
      RECT 296.97 0.18 297.23 8.7 ;
      RECT 297.48 0.17 298.25 0.43 ;
      RECT 297.48 0.17 297.74 8.7 ;
      RECT 297.99 0.17 298.25 8.7 ;
      RECT 298.5 0.18 299.27 0.88 ;
      RECT 298.5 0.18 298.76 8.7 ;
      RECT 299.01 0.18 299.27 8.7 ;
      RECT 299.52 0.17 300.29 0.43 ;
      RECT 299.52 0.17 299.78 8.7 ;
      RECT 300.03 0.17 300.29 8.7 ;
      RECT 300.54 0.18 301.31 0.88 ;
      RECT 300.54 0.18 300.8 8.7 ;
      RECT 301.05 0.18 301.31 8.7 ;
      RECT 284.425 384.61 284.785 385.34 ;
      RECT 284.995 384.61 285.195 385.34 ;
      RECT 302.935 0.18 303.705 0.88 ;
      RECT 302.935 0.18 303.195 8.7 ;
      RECT 303.445 0.18 303.705 8.7 ;
      RECT 303.955 0.17 304.725 0.43 ;
      RECT 303.955 0.17 304.215 8.7 ;
      RECT 304.465 0.17 304.725 8.7 ;
      RECT 285.82 384.53 286.02 385.34 ;
      RECT 301.915 0.3 302.175 8.7 ;
      RECT 305.995 0.18 306.765 0.88 ;
      RECT 305.995 0.18 306.255 8.7 ;
      RECT 306.505 0.18 306.765 8.7 ;
      RECT 302.425 0.3 302.685 8.7 ;
      RECT 304.975 0 305.235 8.7 ;
      RECT 305.485 0 305.745 8.7 ;
      RECT 307.015 0.52 307.275 8.7 ;
      RECT 307.525 0.3 307.785 8.7 ;
      RECT 308.035 0.3 308.295 8.7 ;
      RECT 308.545 0.3 308.805 8.7 ;
      RECT 309.055 0.3 309.315 8.7 ;
      RECT 309.565 0.3 309.825 8.7 ;
      RECT 310.075 0.3 310.335 8.7 ;
      RECT 310.585 0.3 310.845 8.7 ;
      RECT 312.625 0.18 313.395 0.88 ;
      RECT 312.625 0.18 312.885 8.7 ;
      RECT 313.135 0.18 313.395 8.7 ;
      RECT 311.095 0.3 311.355 8.7 ;
      RECT 311.605 0.52 311.865 8.7 ;
      RECT 312.115 0.52 312.375 8.7 ;
      RECT 313.645 0.52 313.905 8.7 ;
      RECT 314.155 0.52 314.415 8.7 ;
      RECT 314.665 0.52 314.925 8.7 ;
      RECT 315.175 0.52 315.435 8.7 ;
      RECT 315.685 0.52 315.945 8.7 ;
      RECT 316.195 0.52 316.455 8.7 ;
      RECT 316.705 0.52 316.965 8.7 ;
      RECT 317.215 0.52 317.475 8.7 ;
      RECT 317.725 0.52 317.985 8.7 ;
      RECT 318.235 0.52 318.495 8.7 ;
      RECT 318.745 0.3 319.005 8.7 ;
      RECT 319.255 0.3 319.515 8.7 ;
      RECT 319.765 0.3 320.025 8.7 ;
      RECT 320.275 0.52 320.535 8.7 ;
      RECT 320.785 0.52 321.045 8.7 ;
      RECT 321.295 0.3 321.555 8.7 ;
      RECT 321.805 0.3 322.065 8.7 ;
      RECT 322.315 0.3 322.575 8.7 ;
      RECT 322.825 0.52 323.085 8.7 ;
      RECT 323.335 0.52 323.595 8.7 ;
      RECT 323.845 0.3 324.105 8.7 ;
      RECT 324.355 0.52 324.615 8.7 ;
      RECT 324.865 0.52 325.125 8.7 ;
      RECT 325.375 0.52 325.635 8.7 ;
      RECT 325.885 0.52 326.145 8.7 ;
      RECT 326.395 0.52 326.655 8.7 ;
      RECT 326.905 0.3 327.165 8.7 ;
      RECT 327.415 0.52 327.675 8.7 ;
      RECT 327.925 0.52 328.185 8.7 ;
      RECT 328.435 0.3 328.695 8.7 ;
      RECT 328.945 0.52 329.205 8.7 ;
      RECT 330.985 0.17 331.755 0.43 ;
      RECT 330.985 0.17 331.245 8.7 ;
      RECT 331.495 0.17 331.755 8.7 ;
      RECT 329.455 0.52 329.715 8.7 ;
      RECT 329.965 0.3 330.225 8.7 ;
      RECT 330.475 0.3 330.735 8.7 ;
      RECT 333.535 0.17 334.305 0.43 ;
      RECT 333.535 0.17 333.795 8.7 ;
      RECT 334.045 0.17 334.305 8.7 ;
      RECT 332.005 0.3 332.265 8.7 ;
      RECT 335.065 0.18 335.835 0.88 ;
      RECT 335.065 0.18 335.325 8.7 ;
      RECT 335.575 0.18 335.835 8.7 ;
      RECT 332.515 0.3 332.775 8.7 ;
      RECT 333.025 0.3 333.285 8.7 ;
      RECT 334.555 0.3 334.815 8.7 ;
      RECT 336.085 0 336.345 8.7 ;
      RECT 336.595 0 336.855 8.7 ;
      RECT 337.105 0.52 337.365 8.7 ;
      RECT 337.615 0.52 337.875 8.7 ;
      RECT 338.125 0.52 338.385 8.7 ;
      RECT 338.635 0.52 338.895 8.7 ;
      RECT 339.145 0 339.405 8.7 ;
      RECT 339.655 0 339.915 8.7 ;
      RECT 340.165 0.3 340.425 8.7 ;
      RECT 340.675 0.3 340.935 8.7 ;
      RECT 341.185 0 341.445 8.7 ;
      RECT 341.695 0 341.955 8.7 ;
      RECT 342.205 0.3 342.465 8.7 ;
      RECT 343.025 0.3 343.285 8.7 ;
      RECT 343.535 0 343.795 8.7 ;
      RECT 344.045 0 344.305 8.7 ;
      RECT 344.555 0.3 344.815 8.7 ;
      RECT 345.065 0.3 345.325 8.7 ;
      RECT 345.575 0 345.835 8.7 ;
      RECT 346.085 0 346.345 8.7 ;
      RECT 346.595 0.52 346.855 8.7 ;
      RECT 347.105 0.52 347.365 8.7 ;
      RECT 347.615 0.52 347.875 8.7 ;
      RECT 349.655 0.18 350.425 0.88 ;
      RECT 349.655 0.18 349.915 8.7 ;
      RECT 350.165 0.18 350.425 8.7 ;
      RECT 348.125 0.52 348.385 8.7 ;
      RECT 351.185 0.17 351.955 0.43 ;
      RECT 351.185 0.17 351.445 8.7 ;
      RECT 351.695 0.17 351.955 8.7 ;
      RECT 348.635 0 348.895 8.7 ;
      RECT 349.145 0 349.405 8.7 ;
      RECT 350.675 0.3 350.935 8.7 ;
      RECT 353.735 0.17 354.505 0.43 ;
      RECT 353.735 0.17 353.995 8.7 ;
      RECT 354.245 0.17 354.505 8.7 ;
      RECT 352.205 0.3 352.465 8.7 ;
      RECT 352.715 0.3 352.975 8.7 ;
      RECT 353.225 0.3 353.485 8.7 ;
      RECT 354.755 0.3 355.015 8.7 ;
      RECT 355.265 0.3 355.525 8.7 ;
      RECT 355.775 0.52 356.035 8.7 ;
      RECT 356.285 0.52 356.545 8.7 ;
      RECT 356.795 0.3 357.055 8.7 ;
      RECT 357.305 0.52 357.565 8.7 ;
      RECT 357.815 0.52 358.075 8.7 ;
      RECT 358.325 0.3 358.585 8.7 ;
      RECT 358.835 0.52 359.095 8.7 ;
      RECT 359.345 0.52 359.605 8.7 ;
      RECT 359.855 0.52 360.115 8.7 ;
      RECT 360.365 0.52 360.625 8.7 ;
      RECT 360.875 0.52 361.135 8.7 ;
      RECT 361.385 0.3 361.645 8.7 ;
      RECT 361.895 0.52 362.155 8.7 ;
      RECT 362.405 0.52 362.665 8.7 ;
      RECT 362.915 0.3 363.175 8.7 ;
      RECT 363.425 0.3 363.685 8.7 ;
      RECT 363.935 0.3 364.195 8.7 ;
      RECT 364.445 0.52 364.705 8.7 ;
      RECT 364.955 0.52 365.215 8.7 ;
      RECT 365.465 0.3 365.725 8.7 ;
      RECT 365.975 0.3 366.235 8.7 ;
      RECT 366.485 0.3 366.745 8.7 ;
      RECT 366.995 0.52 367.255 8.7 ;
      RECT 367.505 0.52 367.765 8.7 ;
      RECT 368.015 0.52 368.275 8.7 ;
      RECT 368.525 0.52 368.785 8.7 ;
      RECT 369.035 0.52 369.295 8.7 ;
      RECT 369.545 0.52 369.805 8.7 ;
      RECT 370.055 0.52 370.315 8.7 ;
      RECT 372.095 0.18 372.865 0.88 ;
      RECT 372.095 0.18 372.355 8.7 ;
      RECT 372.605 0.18 372.865 8.7 ;
      RECT 370.565 0.52 370.825 8.7 ;
      RECT 371.075 0.52 371.335 8.7 ;
      RECT 371.585 0.52 371.845 8.7 ;
      RECT 373.115 0.52 373.375 8.7 ;
      RECT 373.625 0.52 373.885 8.7 ;
      RECT 374.135 0.3 374.395 8.7 ;
      RECT 374.645 0.3 374.905 8.7 ;
      RECT 375.155 0.3 375.415 8.7 ;
      RECT 375.665 0.3 375.925 8.7 ;
      RECT 376.175 0.3 376.435 8.7 ;
      RECT 376.685 0.3 376.945 8.7 ;
      RECT 378.725 0.18 379.495 0.88 ;
      RECT 378.725 0.18 378.985 8.7 ;
      RECT 379.235 0.18 379.495 8.7 ;
      RECT 377.195 0.3 377.455 8.7 ;
      RECT 377.705 0.3 377.965 8.7 ;
      RECT 380.765 0.17 381.535 0.43 ;
      RECT 380.765 0.17 381.025 8.7 ;
      RECT 381.275 0.17 381.535 8.7 ;
      RECT 381.785 0.18 382.555 0.88 ;
      RECT 381.785 0.18 382.045 8.7 ;
      RECT 382.295 0.18 382.555 8.7 ;
      RECT 378.215 0.52 378.475 8.7 ;
      RECT 379.745 0 380.005 8.7 ;
      RECT 384.18 0.18 384.95 0.88 ;
      RECT 384.18 0.18 384.44 8.7 ;
      RECT 384.69 0.18 384.95 8.7 ;
      RECT 385.2 0.17 385.97 0.43 ;
      RECT 385.2 0.17 385.46 8.7 ;
      RECT 385.71 0.17 385.97 8.7 ;
      RECT 386.22 0.18 386.99 0.88 ;
      RECT 386.22 0.18 386.48 8.7 ;
      RECT 386.73 0.18 386.99 8.7 ;
      RECT 387.24 0.17 388.01 0.43 ;
      RECT 387.24 0.17 387.5 8.7 ;
      RECT 387.75 0.17 388.01 8.7 ;
      RECT 388.26 0.18 389.03 0.88 ;
      RECT 388.26 0.18 388.52 8.7 ;
      RECT 388.77 0.18 389.03 8.7 ;
      RECT 389.28 0.17 390.05 0.43 ;
      RECT 389.28 0.17 389.54 8.7 ;
      RECT 389.79 0.17 390.05 8.7 ;
      RECT 390.3 0.18 391.07 0.88 ;
      RECT 390.3 0.18 390.56 8.7 ;
      RECT 390.81 0.18 391.07 8.7 ;
      RECT 391.32 0.17 392.09 0.43 ;
      RECT 391.32 0.17 391.58 8.7 ;
      RECT 391.83 0.17 392.09 8.7 ;
      RECT 392.34 0.18 393.11 0.88 ;
      RECT 392.34 0.18 392.6 8.7 ;
      RECT 392.85 0.18 393.11 8.7 ;
      RECT 393.36 0.17 394.13 0.43 ;
      RECT 393.36 0.17 393.62 8.7 ;
      RECT 393.87 0.17 394.13 8.7 ;
      RECT 394.38 0.18 395.15 0.88 ;
      RECT 394.38 0.18 394.64 8.7 ;
      RECT 394.89 0.18 395.15 8.7 ;
      RECT 395.4 0.17 396.17 0.43 ;
      RECT 395.4 0.17 395.66 8.7 ;
      RECT 395.91 0.17 396.17 8.7 ;
      RECT 396.42 0.18 397.19 0.88 ;
      RECT 396.42 0.18 396.68 8.7 ;
      RECT 396.93 0.18 397.19 8.7 ;
      RECT 397.44 0.17 398.21 0.43 ;
      RECT 397.44 0.17 397.7 8.7 ;
      RECT 397.95 0.17 398.21 8.7 ;
      RECT 398.46 0.18 399.23 0.88 ;
      RECT 398.46 0.18 398.72 8.7 ;
      RECT 398.97 0.18 399.23 8.7 ;
      RECT 380.255 0 380.515 8.7 ;
      RECT 399.48 0.17 400.25 0.43 ;
      RECT 399.48 0.17 399.74 8.7 ;
      RECT 399.99 0.17 400.25 8.7 ;
      RECT 382.805 0.3 383.065 8.7 ;
      RECT 383.315 0.3 383.575 8.7 ;
      RECT 399.47 384.53 399.67 385.34 ;
      RECT 400.295 384.61 400.495 385.34 ;
      RECT 400.705 384.61 401.065 385.34 ;
      RECT 401.01 0.52 401.27 4.315 ;
      RECT 401.275 384.61 401.475 385.34 ;
      RECT 401.93 384.61 402.13 385.34 ;
      RECT 402.185 0.52 402.445 2.82 ;
      RECT 402.34 384.61 402.7 385.34 ;
      RECT 402.995 384.61 403.195 385.34 ;
      RECT 403.49 384.61 403.85 385.34 ;
      RECT 404.425 0.18 405.195 0.88 ;
      RECT 404.425 0.18 404.685 12.9 ;
      RECT 404.935 0.18 405.195 12.9 ;
      RECT 403.715 0.52 403.975 2.82 ;
      RECT 404.06 384.61 404.26 385.34 ;
      RECT 405.445 0.155 406.215 0.445 ;
      RECT 405.445 0.155 405.705 13.21 ;
      RECT 405.955 0.155 406.215 13.21 ;
      RECT 404.715 384.61 404.915 385.34 ;
      RECT 405.125 384.61 405.485 385.34 ;
      RECT 405.695 384.61 405.895 385.34 ;
      RECT 406.35 384.61 406.55 385.34 ;
      RECT 406.76 384.61 407.12 385.34 ;
      RECT 407.415 384.61 407.615 385.34 ;
      RECT 407.91 384.61 408.27 385.34 ;
      RECT 408.15 0.52 408.41 14.115 ;
      RECT 408.48 384.61 408.68 385.34 ;
      RECT 408.66 0.52 408.92 13.45 ;
      RECT 409.135 384.61 409.335 385.34 ;
      RECT 409.68 0.155 410.45 0.445 ;
      RECT 409.68 0.155 409.94 8.665 ;
      RECT 410.19 0.155 410.45 8.665 ;
      RECT 409.17 0.52 409.43 11.315 ;
      RECT 409.545 384.61 409.905 385.34 ;
      RECT 410.115 384.61 410.315 385.34 ;
      RECT 410.7 0.52 410.96 9.955 ;
      RECT 410.77 384.61 410.97 385.34 ;
      RECT 411.18 384.61 411.54 385.34 ;
      RECT 411.835 384.61 412.035 385.34 ;
      RECT 412.33 384.61 412.69 385.34 ;
      RECT 412.74 0.3 413 8.7 ;
      RECT 412.9 384.61 413.1 385.34 ;
      RECT 413.555 384.61 413.755 385.34 ;
      RECT 413.25 0.18 414.02 0.88 ;
      RECT 413.965 384.61 414.325 385.34 ;
      RECT 414.535 384.61 414.735 385.34 ;
      RECT 415.19 384.61 415.39 385.34 ;
      RECT 415.445 0.52 415.705 6.28 ;
      RECT 415.6 384.61 415.96 385.34 ;
      RECT 416.255 384.61 416.455 385.34 ;
      RECT 416.82 0.52 417.08 5.57 ;
      RECT 416.75 384.61 417.11 385.34 ;
      RECT 417.32 384.61 417.52 385.34 ;
      RECT 417.33 0.3 417.59 5.235 ;
      RECT 417.84 0.52 418.1 7.78 ;
      RECT 417.975 384.61 418.175 385.34 ;
      RECT 418.385 384.61 418.745 385.34 ;
      RECT 418.69 0.52 418.95 4.315 ;
      RECT 418.955 384.61 419.155 385.34 ;
      RECT 419.61 384.61 419.81 385.34 ;
      RECT 419.865 0.52 420.125 2.82 ;
      RECT 420.02 384.61 420.38 385.34 ;
      RECT 420.675 384.61 420.875 385.34 ;
      RECT 421.17 384.61 421.53 385.34 ;
      RECT 422.105 0.18 422.875 0.88 ;
      RECT 422.105 0.18 422.365 12.9 ;
      RECT 422.615 0.18 422.875 12.9 ;
      RECT 421.395 0.52 421.655 2.82 ;
      RECT 421.74 384.61 421.94 385.34 ;
      RECT 423.125 0.155 423.895 0.445 ;
      RECT 423.125 0.155 423.385 13.21 ;
      RECT 423.635 0.155 423.895 13.21 ;
      RECT 422.395 384.61 422.595 385.34 ;
      RECT 422.805 384.61 423.165 385.34 ;
      RECT 423.375 384.61 423.575 385.34 ;
      RECT 424.03 384.61 424.23 385.34 ;
      RECT 424.44 384.61 424.8 385.34 ;
      RECT 425.095 384.61 425.295 385.34 ;
      RECT 425.59 384.61 425.95 385.34 ;
      RECT 425.83 0.52 426.09 14.115 ;
      RECT 426.16 384.61 426.36 385.34 ;
      RECT 426.34 0.52 426.6 13.45 ;
      RECT 426.815 384.61 427.015 385.34 ;
      RECT 427.36 0.155 428.13 0.445 ;
      RECT 427.36 0.155 427.62 8.665 ;
      RECT 427.87 0.155 428.13 8.665 ;
      RECT 426.85 0.52 427.11 11.315 ;
      RECT 427.225 384.61 427.585 385.34 ;
      RECT 427.795 384.61 427.995 385.34 ;
      RECT 428.38 0.52 428.64 9.955 ;
      RECT 428.45 384.61 428.65 385.34 ;
      RECT 428.86 384.61 429.22 385.34 ;
      RECT 429.515 384.61 429.715 385.34 ;
      RECT 430.01 384.61 430.37 385.34 ;
      RECT 430.42 0.3 430.68 8.7 ;
      RECT 430.58 384.61 430.78 385.34 ;
      RECT 431.235 384.61 431.435 385.34 ;
      RECT 430.93 0.18 431.7 0.88 ;
      RECT 431.645 384.61 432.005 385.34 ;
      RECT 432.215 384.61 432.415 385.34 ;
      RECT 432.87 384.61 433.07 385.34 ;
      RECT 433.125 0.52 433.385 6.28 ;
      RECT 433.28 384.61 433.64 385.34 ;
      RECT 433.935 384.61 434.135 385.34 ;
      RECT 434.5 0.52 434.76 5.57 ;
      RECT 434.43 384.61 434.79 385.34 ;
      RECT 435 384.61 435.2 385.34 ;
      RECT 435.01 0.3 435.27 5.235 ;
      RECT 435.52 0.52 435.78 7.78 ;
      RECT 435.655 384.61 435.855 385.34 ;
      RECT 436.065 384.61 436.425 385.34 ;
      RECT 436.37 0.52 436.63 4.315 ;
      RECT 436.635 384.61 436.835 385.34 ;
      RECT 437.29 384.61 437.49 385.34 ;
      RECT 437.545 0.52 437.805 2.82 ;
      RECT 437.7 384.61 438.06 385.34 ;
      RECT 438.355 384.61 438.555 385.34 ;
      RECT 438.85 384.61 439.21 385.34 ;
      RECT 439.785 0.18 440.555 0.88 ;
      RECT 439.785 0.18 440.045 12.9 ;
      RECT 440.295 0.18 440.555 12.9 ;
      RECT 439.075 0.52 439.335 2.82 ;
      RECT 439.42 384.61 439.62 385.34 ;
      RECT 440.805 0.155 441.575 0.445 ;
      RECT 440.805 0.155 441.065 13.21 ;
      RECT 441.315 0.155 441.575 13.21 ;
      RECT 440.075 384.61 440.275 385.34 ;
      RECT 440.485 384.61 440.845 385.34 ;
      RECT 441.055 384.61 441.255 385.34 ;
      RECT 441.71 384.61 441.91 385.34 ;
      RECT 442.12 384.61 442.48 385.34 ;
      RECT 442.775 384.61 442.975 385.34 ;
      RECT 443.27 384.61 443.63 385.34 ;
      RECT 443.51 0.52 443.77 14.115 ;
      RECT 443.84 384.61 444.04 385.34 ;
      RECT 444.02 0.52 444.28 13.45 ;
      RECT 444.495 384.61 444.695 385.34 ;
      RECT 445.04 0.155 445.81 0.445 ;
      RECT 445.04 0.155 445.3 8.665 ;
      RECT 445.55 0.155 445.81 8.665 ;
      RECT 444.53 0.52 444.79 11.315 ;
      RECT 444.905 384.61 445.265 385.34 ;
      RECT 445.475 384.61 445.675 385.34 ;
      RECT 446.06 0.52 446.32 9.955 ;
      RECT 446.13 384.61 446.33 385.34 ;
      RECT 446.54 384.61 446.9 385.34 ;
      RECT 447.195 384.61 447.395 385.34 ;
      RECT 447.69 384.61 448.05 385.34 ;
      RECT 448.1 0.3 448.36 8.7 ;
      RECT 448.26 384.61 448.46 385.34 ;
      RECT 448.915 384.61 449.115 385.34 ;
      RECT 448.61 0.18 449.38 0.88 ;
      RECT 449.325 384.61 449.685 385.34 ;
      RECT 449.895 384.61 450.095 385.34 ;
      RECT 450.55 384.61 450.75 385.34 ;
      RECT 450.805 0.52 451.065 6.28 ;
      RECT 450.96 384.61 451.32 385.34 ;
      RECT 451.615 384.61 451.815 385.34 ;
      RECT 452.18 0.52 452.44 5.57 ;
      RECT 452.11 384.61 452.47 385.34 ;
      RECT 452.68 384.61 452.88 385.34 ;
      RECT 452.69 0.3 452.95 5.235 ;
      RECT 453.2 0.52 453.46 7.78 ;
      RECT 453.335 384.61 453.535 385.34 ;
      RECT 453.745 384.61 454.105 385.34 ;
      RECT 454.05 0.52 454.31 4.315 ;
      RECT 454.315 384.61 454.515 385.34 ;
      RECT 454.97 384.61 455.17 385.34 ;
      RECT 455.225 0.52 455.485 2.82 ;
      RECT 455.38 384.61 455.74 385.34 ;
      RECT 456.035 384.61 456.235 385.34 ;
      RECT 456.53 384.61 456.89 385.34 ;
      RECT 457.465 0.18 458.235 0.88 ;
      RECT 457.465 0.18 457.725 12.9 ;
      RECT 457.975 0.18 458.235 12.9 ;
      RECT 456.755 0.52 457.015 2.82 ;
      RECT 457.1 384.61 457.3 385.34 ;
      RECT 458.485 0.155 459.255 0.445 ;
      RECT 458.485 0.155 458.745 13.21 ;
      RECT 458.995 0.155 459.255 13.21 ;
      RECT 457.755 384.61 457.955 385.34 ;
      RECT 458.165 384.61 458.525 385.34 ;
      RECT 458.735 384.61 458.935 385.34 ;
      RECT 459.39 384.61 459.59 385.34 ;
      RECT 459.8 384.61 460.16 385.34 ;
      RECT 460.455 384.61 460.655 385.34 ;
      RECT 460.95 384.61 461.31 385.34 ;
      RECT 461.19 0.52 461.45 14.115 ;
      RECT 461.52 384.61 461.72 385.34 ;
      RECT 461.7 0.52 461.96 13.45 ;
      RECT 462.175 384.61 462.375 385.34 ;
      RECT 462.72 0.155 463.49 0.445 ;
      RECT 462.72 0.155 462.98 8.665 ;
      RECT 463.23 0.155 463.49 8.665 ;
      RECT 462.21 0.52 462.47 11.315 ;
      RECT 462.585 384.61 462.945 385.34 ;
      RECT 463.155 384.61 463.355 385.34 ;
      RECT 463.74 0.52 464 9.955 ;
      RECT 463.81 384.61 464.01 385.34 ;
      RECT 464.22 384.61 464.58 385.34 ;
      RECT 464.875 384.61 465.075 385.34 ;
      RECT 465.37 384.61 465.73 385.34 ;
      RECT 465.78 0.3 466.04 8.7 ;
      RECT 465.94 384.61 466.14 385.34 ;
      RECT 466.595 384.61 466.795 385.34 ;
      RECT 466.29 0.18 467.06 0.88 ;
      RECT 467.005 384.61 467.365 385.34 ;
      RECT 467.575 384.61 467.775 385.34 ;
      RECT 468.23 384.61 468.43 385.34 ;
      RECT 468.485 0.52 468.745 6.28 ;
      RECT 468.64 384.61 469 385.34 ;
      RECT 469.295 384.61 469.495 385.34 ;
      RECT 469.86 0.52 470.12 5.57 ;
      RECT 469.79 384.61 470.15 385.34 ;
      RECT 470.36 384.61 470.56 385.34 ;
      RECT 470.37 0.3 470.63 5.235 ;
      RECT 470.88 0.52 471.14 7.78 ;
      RECT 471.015 384.61 471.215 385.34 ;
      RECT 471.425 384.61 471.785 385.34 ;
      RECT 471.73 0.52 471.99 4.315 ;
      RECT 471.995 384.61 472.195 385.34 ;
      RECT 472.65 384.61 472.85 385.34 ;
      RECT 472.905 0.52 473.165 2.82 ;
      RECT 473.06 384.61 473.42 385.34 ;
      RECT 473.715 384.61 473.915 385.34 ;
      RECT 474.21 384.61 474.57 385.34 ;
      RECT 475.145 0.18 475.915 0.88 ;
      RECT 475.145 0.18 475.405 12.9 ;
      RECT 475.655 0.18 475.915 12.9 ;
      RECT 474.435 0.52 474.695 2.82 ;
      RECT 474.78 384.61 474.98 385.34 ;
      RECT 476.165 0.155 476.935 0.445 ;
      RECT 476.165 0.155 476.425 13.21 ;
      RECT 476.675 0.155 476.935 13.21 ;
      RECT 475.435 384.61 475.635 385.34 ;
      RECT 475.845 384.61 476.205 385.34 ;
      RECT 476.415 384.61 476.615 385.34 ;
      RECT 477.07 384.61 477.27 385.34 ;
      RECT 477.48 384.61 477.84 385.34 ;
      RECT 478.135 384.61 478.335 385.34 ;
      RECT 478.63 384.61 478.99 385.34 ;
      RECT 478.87 0.52 479.13 14.115 ;
      RECT 479.2 384.61 479.4 385.34 ;
      RECT 479.38 0.52 479.64 13.45 ;
      RECT 479.855 384.61 480.055 385.34 ;
      RECT 480.4 0.155 481.17 0.445 ;
      RECT 480.4 0.155 480.66 8.665 ;
      RECT 480.91 0.155 481.17 8.665 ;
      RECT 479.89 0.52 480.15 11.315 ;
      RECT 480.265 384.61 480.625 385.34 ;
      RECT 480.835 384.61 481.035 385.34 ;
      RECT 481.42 0.52 481.68 9.955 ;
      RECT 481.49 384.61 481.69 385.34 ;
      RECT 481.9 384.61 482.26 385.34 ;
      RECT 482.555 384.61 482.755 385.34 ;
      RECT 483.05 384.61 483.41 385.34 ;
      RECT 483.46 0.3 483.72 8.7 ;
      RECT 483.62 384.61 483.82 385.34 ;
      RECT 484.275 384.61 484.475 385.34 ;
      RECT 483.97 0.18 484.74 0.88 ;
      RECT 484.685 384.61 485.045 385.34 ;
      RECT 485.255 384.61 485.455 385.34 ;
      RECT 485.91 384.61 486.11 385.34 ;
      RECT 486.165 0.52 486.425 6.28 ;
      RECT 486.32 384.61 486.68 385.34 ;
      RECT 486.975 384.61 487.175 385.34 ;
      RECT 487.54 0.52 487.8 5.57 ;
      RECT 487.47 384.61 487.83 385.34 ;
      RECT 488.04 384.61 488.24 385.34 ;
      RECT 488.05 0.3 488.31 5.235 ;
      RECT 488.56 0.52 488.82 7.78 ;
      RECT 488.695 384.61 488.895 385.34 ;
      RECT 489.105 384.61 489.465 385.34 ;
      RECT 489.41 0.52 489.67 4.315 ;
      RECT 489.675 384.61 489.875 385.34 ;
      RECT 490.33 384.61 490.53 385.34 ;
      RECT 490.585 0.52 490.845 2.82 ;
      RECT 490.74 384.61 491.1 385.34 ;
      RECT 491.395 384.61 491.595 385.34 ;
      RECT 491.89 384.61 492.25 385.34 ;
      RECT 492.825 0.18 493.595 0.88 ;
      RECT 492.825 0.18 493.085 12.9 ;
      RECT 493.335 0.18 493.595 12.9 ;
      RECT 492.115 0.52 492.375 2.82 ;
      RECT 492.46 384.61 492.66 385.34 ;
      RECT 493.845 0.155 494.615 0.445 ;
      RECT 493.845 0.155 494.105 13.21 ;
      RECT 494.355 0.155 494.615 13.21 ;
      RECT 493.115 384.61 493.315 385.34 ;
      RECT 493.525 384.61 493.885 385.34 ;
      RECT 494.095 384.61 494.295 385.34 ;
      RECT 494.75 384.61 494.95 385.34 ;
      RECT 495.16 384.61 495.52 385.34 ;
      RECT 495.815 384.61 496.015 385.34 ;
      RECT 496.31 384.61 496.67 385.34 ;
      RECT 496.55 0.52 496.81 14.115 ;
      RECT 496.88 384.61 497.08 385.34 ;
      RECT 497.06 0.52 497.32 13.45 ;
      RECT 497.535 384.61 497.735 385.34 ;
      RECT 498.08 0.155 498.85 0.445 ;
      RECT 498.08 0.155 498.34 8.665 ;
      RECT 498.59 0.155 498.85 8.665 ;
      RECT 497.57 0.52 497.83 11.315 ;
      RECT 497.945 384.61 498.305 385.34 ;
      RECT 498.515 384.61 498.715 385.34 ;
      RECT 499.1 0.52 499.36 9.955 ;
      RECT 499.17 384.61 499.37 385.34 ;
      RECT 499.58 384.61 499.94 385.34 ;
      RECT 500.235 384.61 500.435 385.34 ;
      RECT 500.73 384.61 501.09 385.34 ;
      RECT 501.14 0.3 501.4 8.7 ;
      RECT 501.3 384.61 501.5 385.34 ;
      RECT 501.955 384.61 502.155 385.34 ;
      RECT 501.65 0.18 502.42 0.88 ;
      RECT 502.365 384.61 502.725 385.34 ;
      RECT 502.935 384.61 503.135 385.34 ;
      RECT 503.59 384.61 503.79 385.34 ;
      RECT 503.845 0.52 504.105 6.28 ;
      RECT 504 384.61 504.36 385.34 ;
      RECT 504.655 384.61 504.855 385.34 ;
      RECT 505.22 0.52 505.48 5.57 ;
      RECT 505.15 384.61 505.51 385.34 ;
      RECT 505.72 384.61 505.92 385.34 ;
      RECT 505.73 0.3 505.99 5.235 ;
      RECT 506.24 0.52 506.5 7.78 ;
      RECT 506.375 384.61 506.575 385.34 ;
      RECT 506.785 384.61 507.145 385.34 ;
      RECT 507.09 0.52 507.35 4.315 ;
      RECT 507.355 384.61 507.555 385.34 ;
      RECT 508.01 384.61 508.21 385.34 ;
      RECT 508.265 0.52 508.525 2.82 ;
      RECT 508.42 384.61 508.78 385.34 ;
      RECT 509.075 384.61 509.275 385.34 ;
      RECT 509.57 384.61 509.93 385.34 ;
      RECT 510.505 0.18 511.275 0.88 ;
      RECT 510.505 0.18 510.765 12.9 ;
      RECT 511.015 0.18 511.275 12.9 ;
      RECT 509.795 0.52 510.055 2.82 ;
      RECT 510.14 384.61 510.34 385.34 ;
      RECT 511.525 0.155 512.295 0.445 ;
      RECT 511.525 0.155 511.785 13.21 ;
      RECT 512.035 0.155 512.295 13.21 ;
      RECT 510.795 384.61 510.995 385.34 ;
      RECT 511.205 384.61 511.565 385.34 ;
      RECT 511.775 384.61 511.975 385.34 ;
      RECT 512.43 384.61 512.63 385.34 ;
      RECT 512.84 384.61 513.2 385.34 ;
      RECT 513.495 384.61 513.695 385.34 ;
      RECT 513.99 384.61 514.35 385.34 ;
      RECT 514.23 0.52 514.49 14.115 ;
      RECT 514.56 384.61 514.76 385.34 ;
      RECT 514.74 0.52 515 13.45 ;
      RECT 515.215 384.61 515.415 385.34 ;
      RECT 515.76 0.155 516.53 0.445 ;
      RECT 515.76 0.155 516.02 8.665 ;
      RECT 516.27 0.155 516.53 8.665 ;
      RECT 515.25 0.52 515.51 11.315 ;
      RECT 515.625 384.61 515.985 385.34 ;
      RECT 516.195 384.61 516.395 385.34 ;
      RECT 516.78 0.52 517.04 9.955 ;
      RECT 516.85 384.61 517.05 385.34 ;
      RECT 517.26 384.61 517.62 385.34 ;
      RECT 517.915 384.61 518.115 385.34 ;
      RECT 518.41 384.61 518.77 385.34 ;
      RECT 518.82 0.3 519.08 8.7 ;
      RECT 518.98 384.61 519.18 385.34 ;
      RECT 519.635 384.61 519.835 385.34 ;
      RECT 519.33 0.18 520.1 0.88 ;
      RECT 520.045 384.61 520.405 385.34 ;
      RECT 520.615 384.61 520.815 385.34 ;
      RECT 521.27 384.61 521.47 385.34 ;
      RECT 521.525 0.52 521.785 6.28 ;
      RECT 521.68 384.61 522.04 385.34 ;
      RECT 522.335 384.61 522.535 385.34 ;
      RECT 522.9 0.52 523.16 5.57 ;
      RECT 522.83 384.61 523.19 385.34 ;
      RECT 523.4 384.61 523.6 385.34 ;
      RECT 523.41 0.3 523.67 5.235 ;
      RECT 523.92 0.52 524.18 7.78 ;
      RECT 524.055 384.61 524.255 385.34 ;
      RECT 524.465 384.61 524.825 385.34 ;
      RECT 524.77 0.52 525.03 4.315 ;
      RECT 525.035 384.61 525.235 385.34 ;
      RECT 525.69 384.61 525.89 385.34 ;
      RECT 525.945 0.52 526.205 2.82 ;
      RECT 526.1 384.61 526.46 385.34 ;
      RECT 526.755 384.61 526.955 385.34 ;
      RECT 527.25 384.61 527.61 385.34 ;
      RECT 528.185 0.18 528.955 0.88 ;
      RECT 528.185 0.18 528.445 12.9 ;
      RECT 528.695 0.18 528.955 12.9 ;
      RECT 527.475 0.52 527.735 2.82 ;
      RECT 527.82 384.61 528.02 385.34 ;
      RECT 529.205 0.155 529.975 0.445 ;
      RECT 529.205 0.155 529.465 13.21 ;
      RECT 529.715 0.155 529.975 13.21 ;
      RECT 528.475 384.61 528.675 385.34 ;
      RECT 528.885 384.61 529.245 385.34 ;
      RECT 529.455 384.61 529.655 385.34 ;
      RECT 530.11 384.61 530.31 385.34 ;
      RECT 530.52 384.61 530.88 385.34 ;
      RECT 531.175 384.61 531.375 385.34 ;
      RECT 531.67 384.61 532.03 385.34 ;
      RECT 531.91 0.52 532.17 14.115 ;
      RECT 532.24 384.61 532.44 385.34 ;
      RECT 532.42 0.52 532.68 13.45 ;
      RECT 532.895 384.61 533.095 385.34 ;
      RECT 533.44 0.155 534.21 0.445 ;
      RECT 533.44 0.155 533.7 8.665 ;
      RECT 533.95 0.155 534.21 8.665 ;
      RECT 532.93 0.52 533.19 11.315 ;
      RECT 533.305 384.61 533.665 385.34 ;
      RECT 533.875 384.61 534.075 385.34 ;
      RECT 534.46 0.52 534.72 9.955 ;
      RECT 534.53 384.61 534.73 385.34 ;
      RECT 534.94 384.61 535.3 385.34 ;
      RECT 535.595 384.61 535.795 385.34 ;
      RECT 536.09 384.61 536.45 385.34 ;
      RECT 536.5 0.3 536.76 8.7 ;
      RECT 536.66 384.61 536.86 385.34 ;
      RECT 537.315 384.61 537.515 385.34 ;
      RECT 537.01 0.18 537.78 0.88 ;
      RECT 537.725 384.61 538.085 385.34 ;
      RECT 538.295 384.61 538.495 385.34 ;
      RECT 538.95 384.61 539.15 385.34 ;
      RECT 539.205 0.52 539.465 6.28 ;
      RECT 539.36 384.61 539.72 385.34 ;
      RECT 540.015 384.61 540.215 385.34 ;
      RECT 540.58 0.52 540.84 5.57 ;
      RECT 540.51 384.61 540.87 385.34 ;
      RECT 541.08 384.61 541.28 385.34 ;
      RECT 541.09 0.3 541.35 5.235 ;
      RECT 541.6 0.52 541.86 7.78 ;
      RECT 541.735 384.61 541.935 385.34 ;
      RECT 542.145 384.61 542.505 385.34 ;
      RECT 542.45 0.52 542.71 4.315 ;
      RECT 542.715 384.61 542.915 385.34 ;
      RECT 543.37 384.61 543.57 385.34 ;
      RECT 543.625 0.52 543.885 2.82 ;
      RECT 543.78 384.61 544.14 385.34 ;
      RECT 544.435 384.61 544.635 385.34 ;
      RECT 544.93 384.61 545.29 385.34 ;
      RECT 545.865 0.18 546.635 0.88 ;
      RECT 545.865 0.18 546.125 12.9 ;
      RECT 546.375 0.18 546.635 12.9 ;
      RECT 545.155 0.52 545.415 2.82 ;
      RECT 545.5 384.61 545.7 385.34 ;
      RECT 546.885 0.155 547.655 0.445 ;
      RECT 546.885 0.155 547.145 13.21 ;
      RECT 547.395 0.155 547.655 13.21 ;
      RECT 546.155 384.61 546.355 385.34 ;
      RECT 546.565 384.61 546.925 385.34 ;
      RECT 547.135 384.61 547.335 385.34 ;
      RECT 547.79 384.61 547.99 385.34 ;
      RECT 548.2 384.61 548.56 385.34 ;
      RECT 548.855 384.61 549.055 385.34 ;
      RECT 549.35 384.61 549.71 385.34 ;
      RECT 549.59 0.52 549.85 14.115 ;
      RECT 549.92 384.61 550.12 385.34 ;
      RECT 550.1 0.52 550.36 13.45 ;
      RECT 550.575 384.61 550.775 385.34 ;
      RECT 551.12 0.155 551.89 0.445 ;
      RECT 551.12 0.155 551.38 8.665 ;
      RECT 551.63 0.155 551.89 8.665 ;
      RECT 550.61 0.52 550.87 11.315 ;
      RECT 550.985 384.61 551.345 385.34 ;
      RECT 551.555 384.61 551.755 385.34 ;
      RECT 552.14 0.52 552.4 9.955 ;
      RECT 552.21 384.61 552.41 385.34 ;
      RECT 552.62 384.61 552.98 385.34 ;
      RECT 553.275 384.61 553.475 385.34 ;
      RECT 553.77 384.61 554.13 385.34 ;
      RECT 554.18 0.3 554.44 8.7 ;
      RECT 554.34 384.61 554.54 385.34 ;
      RECT 554.995 384.61 555.195 385.34 ;
      RECT 554.69 0.18 555.46 0.88 ;
      RECT 555.405 384.61 555.765 385.34 ;
      RECT 555.975 384.61 556.175 385.34 ;
      RECT 556.63 384.61 556.83 385.34 ;
      RECT 556.885 0.52 557.145 6.28 ;
      RECT 557.04 384.61 557.4 385.34 ;
      RECT 557.695 384.61 557.895 385.34 ;
      RECT 558.26 0.52 558.52 5.57 ;
      RECT 558.19 384.61 558.55 385.34 ;
      RECT 558.76 384.61 558.96 385.34 ;
      RECT 558.77 0.3 559.03 5.235 ;
      RECT 559.28 0.52 559.54 7.78 ;
      RECT 559.415 384.61 559.615 385.34 ;
      RECT 559.825 384.61 560.185 385.34 ;
      RECT 560.13 0.52 560.39 4.315 ;
      RECT 560.395 384.61 560.595 385.34 ;
      RECT 561.05 384.61 561.25 385.34 ;
      RECT 561.305 0.52 561.565 2.82 ;
      RECT 561.46 384.61 561.82 385.34 ;
      RECT 562.115 384.61 562.315 385.34 ;
      RECT 562.61 384.61 562.97 385.34 ;
      RECT 563.545 0.18 564.315 0.88 ;
      RECT 563.545 0.18 563.805 12.9 ;
      RECT 564.055 0.18 564.315 12.9 ;
      RECT 562.835 0.52 563.095 2.82 ;
      RECT 563.18 384.61 563.38 385.34 ;
      RECT 564.565 0.155 565.335 0.445 ;
      RECT 564.565 0.155 564.825 13.21 ;
      RECT 565.075 0.155 565.335 13.21 ;
      RECT 563.835 384.61 564.035 385.34 ;
      RECT 564.245 384.61 564.605 385.34 ;
      RECT 564.815 384.61 565.015 385.34 ;
      RECT 565.47 384.61 565.67 385.34 ;
      RECT 565.88 384.61 566.24 385.34 ;
      RECT 566.535 384.61 566.735 385.34 ;
      RECT 567.03 384.61 567.39 385.34 ;
      RECT 567.27 0.52 567.53 14.115 ;
      RECT 567.6 384.61 567.8 385.34 ;
      RECT 567.78 0.52 568.04 13.45 ;
      RECT 568.255 384.61 568.455 385.34 ;
      RECT 568.8 0.155 569.57 0.445 ;
      RECT 568.8 0.155 569.06 8.665 ;
      RECT 569.31 0.155 569.57 8.665 ;
      RECT 568.29 0.52 568.55 11.315 ;
      RECT 568.665 384.61 569.025 385.34 ;
      RECT 569.235 384.61 569.435 385.34 ;
      RECT 569.82 0.52 570.08 9.955 ;
      RECT 569.89 384.61 570.09 385.34 ;
      RECT 570.3 384.61 570.66 385.34 ;
      RECT 570.955 384.61 571.155 385.34 ;
      RECT 571.45 384.61 571.81 385.34 ;
      RECT 571.86 0.3 572.12 8.7 ;
      RECT 572.02 384.61 572.22 385.34 ;
      RECT 572.675 384.61 572.875 385.34 ;
      RECT 572.37 0.18 573.14 0.88 ;
      RECT 573.085 384.61 573.445 385.34 ;
      RECT 573.655 384.61 573.855 385.34 ;
      RECT 574.31 384.61 574.51 385.34 ;
      RECT 574.565 0.52 574.825 6.28 ;
      RECT 574.72 384.61 575.08 385.34 ;
      RECT 575.375 384.61 575.575 385.34 ;
      RECT 575.94 0.52 576.2 5.57 ;
      RECT 575.87 384.61 576.23 385.34 ;
      RECT 576.44 384.61 576.64 385.34 ;
      RECT 576.45 0.3 576.71 5.235 ;
      RECT 576.96 0.52 577.22 7.78 ;
      RECT 577.095 384.61 577.295 385.34 ;
      RECT 577.505 384.61 577.865 385.34 ;
      RECT 577.81 0.52 578.07 4.315 ;
      RECT 578.075 384.61 578.275 385.34 ;
      RECT 578.73 384.61 578.93 385.34 ;
      RECT 578.985 0.52 579.245 2.82 ;
      RECT 579.14 384.61 579.5 385.34 ;
      RECT 579.795 384.61 579.995 385.34 ;
      RECT 580.29 384.61 580.65 385.34 ;
      RECT 581.225 0.18 581.995 0.88 ;
      RECT 581.225 0.18 581.485 12.9 ;
      RECT 581.735 0.18 581.995 12.9 ;
      RECT 580.515 0.52 580.775 2.82 ;
      RECT 580.86 384.61 581.06 385.34 ;
      RECT 582.245 0.155 583.015 0.445 ;
      RECT 582.245 0.155 582.505 13.21 ;
      RECT 582.755 0.155 583.015 13.21 ;
      RECT 581.515 384.61 581.715 385.34 ;
      RECT 581.925 384.61 582.285 385.34 ;
      RECT 582.495 384.61 582.695 385.34 ;
      RECT 583.15 384.61 583.35 385.34 ;
      RECT 583.56 384.61 583.92 385.34 ;
      RECT 584.215 384.61 584.415 385.34 ;
      RECT 584.71 384.61 585.07 385.34 ;
      RECT 584.95 0.52 585.21 14.115 ;
      RECT 585.28 384.61 585.48 385.34 ;
      RECT 585.46 0.52 585.72 13.45 ;
      RECT 585.935 384.61 586.135 385.34 ;
      RECT 586.48 0.155 587.25 0.445 ;
      RECT 586.48 0.155 586.74 8.665 ;
      RECT 586.99 0.155 587.25 8.665 ;
      RECT 585.97 0.52 586.23 11.315 ;
      RECT 586.345 384.61 586.705 385.34 ;
      RECT 586.915 384.61 587.115 385.34 ;
      RECT 587.5 0.52 587.76 9.955 ;
      RECT 587.57 384.61 587.77 385.34 ;
      RECT 587.98 384.61 588.34 385.34 ;
      RECT 588.635 384.61 588.835 385.34 ;
      RECT 589.13 384.61 589.49 385.34 ;
      RECT 589.54 0.3 589.8 8.7 ;
      RECT 589.7 384.61 589.9 385.34 ;
      RECT 590.355 384.61 590.555 385.34 ;
      RECT 590.05 0.18 590.82 0.88 ;
      RECT 590.765 384.61 591.125 385.34 ;
      RECT 591.335 384.61 591.535 385.34 ;
      RECT 591.99 384.61 592.19 385.34 ;
      RECT 592.245 0.52 592.505 6.28 ;
      RECT 592.4 384.61 592.76 385.34 ;
      RECT 593.055 384.61 593.255 385.34 ;
      RECT 593.62 0.52 593.88 5.57 ;
      RECT 593.55 384.61 593.91 385.34 ;
      RECT 594.12 384.61 594.32 385.34 ;
      RECT 594.13 0.3 594.39 5.235 ;
      RECT 594.64 0.52 594.9 7.78 ;
      RECT 594.775 384.61 594.975 385.34 ;
      RECT 595.185 384.61 595.545 385.34 ;
      RECT 595.49 0.52 595.75 4.315 ;
      RECT 595.755 384.61 595.955 385.34 ;
      RECT 596.41 384.61 596.61 385.34 ;
      RECT 596.665 0.52 596.925 2.82 ;
      RECT 596.82 384.61 597.18 385.34 ;
      RECT 597.475 384.61 597.675 385.34 ;
      RECT 597.97 384.61 598.33 385.34 ;
      RECT 598.905 0.18 599.675 0.88 ;
      RECT 598.905 0.18 599.165 12.9 ;
      RECT 599.415 0.18 599.675 12.9 ;
      RECT 598.195 0.52 598.455 2.82 ;
      RECT 598.54 384.61 598.74 385.34 ;
      RECT 599.925 0.155 600.695 0.445 ;
      RECT 599.925 0.155 600.185 13.21 ;
      RECT 600.435 0.155 600.695 13.21 ;
      RECT 599.195 384.61 599.395 385.34 ;
      RECT 599.605 384.61 599.965 385.34 ;
      RECT 600.175 384.61 600.375 385.34 ;
      RECT 600.83 384.61 601.03 385.34 ;
      RECT 601.24 384.61 601.6 385.34 ;
      RECT 601.895 384.61 602.095 385.34 ;
      RECT 602.39 384.61 602.75 385.34 ;
      RECT 602.63 0.52 602.89 14.115 ;
      RECT 602.96 384.61 603.16 385.34 ;
      RECT 603.14 0.52 603.4 13.45 ;
      RECT 603.615 384.61 603.815 385.34 ;
      RECT 604.16 0.155 604.93 0.445 ;
      RECT 604.16 0.155 604.42 8.665 ;
      RECT 604.67 0.155 604.93 8.665 ;
      RECT 603.65 0.52 603.91 11.315 ;
      RECT 604.025 384.61 604.385 385.34 ;
      RECT 604.595 384.61 604.795 385.34 ;
      RECT 605.18 0.52 605.44 9.955 ;
      RECT 605.25 384.61 605.45 385.34 ;
      RECT 605.66 384.61 606.02 385.34 ;
      RECT 606.315 384.61 606.515 385.34 ;
      RECT 606.81 384.61 607.17 385.34 ;
      RECT 607.22 0.3 607.48 8.7 ;
      RECT 607.38 384.61 607.58 385.34 ;
      RECT 608.035 384.61 608.235 385.34 ;
      RECT 607.73 0.18 608.5 0.88 ;
      RECT 608.445 384.61 608.805 385.34 ;
      RECT 609.015 384.61 609.215 385.34 ;
      RECT 609.67 384.61 609.87 385.34 ;
      RECT 609.925 0.52 610.185 6.28 ;
      RECT 610.08 384.61 610.44 385.34 ;
      RECT 610.735 384.61 610.935 385.34 ;
      RECT 611.3 0.52 611.56 5.57 ;
      RECT 611.23 384.61 611.59 385.34 ;
      RECT 611.8 384.61 612 385.34 ;
      RECT 611.81 0.3 612.07 5.235 ;
      RECT 612.32 0.52 612.58 7.78 ;
      RECT 612.455 384.61 612.655 385.34 ;
      RECT 612.865 384.61 613.225 385.34 ;
      RECT 613.17 0.52 613.43 4.315 ;
      RECT 613.435 384.61 613.635 385.34 ;
      RECT 614.09 384.61 614.29 385.34 ;
      RECT 614.345 0.52 614.605 2.82 ;
      RECT 614.5 384.61 614.86 385.34 ;
      RECT 615.155 384.61 615.355 385.34 ;
      RECT 615.65 384.61 616.01 385.34 ;
      RECT 616.585 0.18 617.355 0.88 ;
      RECT 616.585 0.18 616.845 12.9 ;
      RECT 617.095 0.18 617.355 12.9 ;
      RECT 615.875 0.52 616.135 2.82 ;
      RECT 616.22 384.61 616.42 385.34 ;
      RECT 617.605 0.155 618.375 0.445 ;
      RECT 617.605 0.155 617.865 13.21 ;
      RECT 618.115 0.155 618.375 13.21 ;
      RECT 616.875 384.61 617.075 385.34 ;
      RECT 617.285 384.61 617.645 385.34 ;
      RECT 617.855 384.61 618.055 385.34 ;
      RECT 618.51 384.61 618.71 385.34 ;
      RECT 618.92 384.61 619.28 385.34 ;
      RECT 619.575 384.61 619.775 385.34 ;
      RECT 620.07 384.61 620.43 385.34 ;
      RECT 620.31 0.52 620.57 14.115 ;
      RECT 620.64 384.61 620.84 385.34 ;
      RECT 620.82 0.52 621.08 13.45 ;
      RECT 621.295 384.61 621.495 385.34 ;
      RECT 621.84 0.155 622.61 0.445 ;
      RECT 621.84 0.155 622.1 8.665 ;
      RECT 622.35 0.155 622.61 8.665 ;
      RECT 621.33 0.52 621.59 11.315 ;
      RECT 621.705 384.61 622.065 385.34 ;
      RECT 622.275 384.61 622.475 385.34 ;
      RECT 622.86 0.52 623.12 9.955 ;
      RECT 622.93 384.61 623.13 385.34 ;
      RECT 623.34 384.61 623.7 385.34 ;
      RECT 623.995 384.61 624.195 385.34 ;
      RECT 624.49 384.61 624.85 385.34 ;
      RECT 624.9 0.3 625.16 8.7 ;
      RECT 625.06 384.61 625.26 385.34 ;
      RECT 625.715 384.61 625.915 385.34 ;
      RECT 625.41 0.18 626.18 0.88 ;
      RECT 626.125 384.61 626.485 385.34 ;
      RECT 626.695 384.61 626.895 385.34 ;
      RECT 627.35 384.61 627.55 385.34 ;
      RECT 627.605 0.52 627.865 6.28 ;
      RECT 627.76 384.61 628.12 385.34 ;
      RECT 628.415 384.61 628.615 385.34 ;
      RECT 628.98 0.52 629.24 5.57 ;
      RECT 628.91 384.61 629.27 385.34 ;
      RECT 629.48 384.61 629.68 385.34 ;
      RECT 629.49 0.3 629.75 5.235 ;
      RECT 630 0.52 630.26 7.78 ;
      RECT 630.135 384.61 630.335 385.34 ;
      RECT 630.545 384.61 630.905 385.34 ;
      RECT 630.85 0.52 631.11 4.315 ;
      RECT 631.115 384.61 631.315 385.34 ;
      RECT 631.77 384.61 631.97 385.34 ;
      RECT 632.025 0.52 632.285 2.82 ;
      RECT 632.18 384.61 632.54 385.34 ;
      RECT 632.835 384.61 633.035 385.34 ;
      RECT 633.33 384.61 633.69 385.34 ;
      RECT 634.265 0.18 635.035 0.88 ;
      RECT 634.265 0.18 634.525 12.9 ;
      RECT 634.775 0.18 635.035 12.9 ;
      RECT 633.555 0.52 633.815 2.82 ;
      RECT 633.9 384.61 634.1 385.34 ;
      RECT 635.285 0.155 636.055 0.445 ;
      RECT 635.285 0.155 635.545 13.21 ;
      RECT 635.795 0.155 636.055 13.21 ;
      RECT 634.555 384.61 634.755 385.34 ;
      RECT 634.965 384.61 635.325 385.34 ;
      RECT 635.535 384.61 635.735 385.34 ;
      RECT 636.19 384.61 636.39 385.34 ;
      RECT 636.6 384.61 636.96 385.34 ;
      RECT 637.255 384.61 637.455 385.34 ;
      RECT 637.75 384.61 638.11 385.34 ;
      RECT 637.99 0.52 638.25 14.115 ;
      RECT 638.32 384.61 638.52 385.34 ;
      RECT 638.5 0.52 638.76 13.45 ;
      RECT 638.975 384.61 639.175 385.34 ;
      RECT 639.52 0.155 640.29 0.445 ;
      RECT 639.52 0.155 639.78 8.665 ;
      RECT 640.03 0.155 640.29 8.665 ;
      RECT 639.01 0.52 639.27 11.315 ;
      RECT 639.385 384.61 639.745 385.34 ;
      RECT 639.955 384.61 640.155 385.34 ;
      RECT 640.54 0.52 640.8 9.955 ;
      RECT 640.61 384.61 640.81 385.34 ;
      RECT 641.02 384.61 641.38 385.34 ;
      RECT 641.675 384.61 641.875 385.34 ;
      RECT 642.17 384.61 642.53 385.34 ;
      RECT 642.58 0.3 642.84 8.7 ;
      RECT 642.74 384.61 642.94 385.34 ;
      RECT 643.395 384.61 643.595 385.34 ;
      RECT 643.09 0.18 643.86 0.88 ;
      RECT 643.805 384.61 644.165 385.34 ;
      RECT 644.375 384.61 644.575 385.34 ;
      RECT 645.03 384.61 645.23 385.34 ;
      RECT 645.285 0.52 645.545 6.28 ;
      RECT 645.44 384.61 645.8 385.34 ;
      RECT 646.095 384.61 646.295 385.34 ;
      RECT 646.66 0.52 646.92 5.57 ;
      RECT 646.59 384.61 646.95 385.34 ;
      RECT 647.16 384.61 647.36 385.34 ;
      RECT 647.17 0.3 647.43 5.235 ;
      RECT 647.68 0.52 647.94 7.78 ;
      RECT 647.815 384.61 648.015 385.34 ;
      RECT 648.225 384.61 648.585 385.34 ;
      RECT 648.53 0.52 648.79 4.315 ;
      RECT 648.795 384.61 648.995 385.34 ;
      RECT 649.45 384.61 649.65 385.34 ;
      RECT 649.705 0.52 649.965 2.82 ;
      RECT 649.86 384.61 650.22 385.34 ;
      RECT 650.515 384.61 650.715 385.34 ;
      RECT 651.01 384.61 651.37 385.34 ;
      RECT 651.945 0.18 652.715 0.88 ;
      RECT 651.945 0.18 652.205 12.9 ;
      RECT 652.455 0.18 652.715 12.9 ;
      RECT 651.235 0.52 651.495 2.82 ;
      RECT 651.58 384.61 651.78 385.34 ;
      RECT 652.965 0.155 653.735 0.445 ;
      RECT 652.965 0.155 653.225 13.21 ;
      RECT 653.475 0.155 653.735 13.21 ;
      RECT 652.235 384.61 652.435 385.34 ;
      RECT 652.645 384.61 653.005 385.34 ;
      RECT 653.215 384.61 653.415 385.34 ;
      RECT 653.87 384.61 654.07 385.34 ;
      RECT 654.28 384.61 654.64 385.34 ;
      RECT 654.935 384.61 655.135 385.34 ;
      RECT 655.43 384.61 655.79 385.34 ;
      RECT 655.67 0.52 655.93 14.115 ;
      RECT 656 384.61 656.2 385.34 ;
      RECT 656.18 0.52 656.44 13.45 ;
      RECT 656.655 384.61 656.855 385.34 ;
      RECT 657.2 0.155 657.97 0.445 ;
      RECT 657.2 0.155 657.46 8.665 ;
      RECT 657.71 0.155 657.97 8.665 ;
      RECT 656.69 0.52 656.95 11.315 ;
      RECT 657.065 384.61 657.425 385.34 ;
      RECT 657.635 384.61 657.835 385.34 ;
      RECT 658.22 0.52 658.48 9.955 ;
      RECT 658.29 384.61 658.49 385.34 ;
      RECT 658.7 384.61 659.06 385.34 ;
      RECT 659.355 384.61 659.555 385.34 ;
      RECT 659.85 384.61 660.21 385.34 ;
      RECT 660.26 0.3 660.52 8.7 ;
      RECT 660.42 384.61 660.62 385.34 ;
      RECT 661.075 384.61 661.275 385.34 ;
      RECT 660.77 0.18 661.54 0.88 ;
      RECT 661.485 384.61 661.845 385.34 ;
      RECT 662.055 384.61 662.255 385.34 ;
      RECT 662.71 384.61 662.91 385.34 ;
      RECT 662.965 0.52 663.225 6.28 ;
      RECT 663.12 384.61 663.48 385.34 ;
      RECT 663.775 384.61 663.975 385.34 ;
      RECT 664.34 0.52 664.6 5.57 ;
      RECT 664.27 384.61 664.63 385.34 ;
      RECT 664.84 384.61 665.04 385.34 ;
      RECT 664.85 0.3 665.11 5.235 ;
      RECT 665.36 0.52 665.62 7.78 ;
      RECT 665.495 384.61 665.695 385.34 ;
      RECT 665.905 384.61 666.265 385.34 ;
      RECT 666.21 0.52 666.47 4.315 ;
      RECT 666.475 384.61 666.675 385.34 ;
      RECT 667.13 384.61 667.33 385.34 ;
      RECT 667.385 0.52 667.645 2.82 ;
      RECT 667.54 384.61 667.9 385.34 ;
      RECT 668.195 384.61 668.395 385.34 ;
      RECT 668.69 384.61 669.05 385.34 ;
      RECT 669.625 0.18 670.395 0.88 ;
      RECT 669.625 0.18 669.885 12.9 ;
      RECT 670.135 0.18 670.395 12.9 ;
      RECT 668.915 0.52 669.175 2.82 ;
      RECT 669.26 384.61 669.46 385.34 ;
      RECT 670.645 0.155 671.415 0.445 ;
      RECT 670.645 0.155 670.905 13.21 ;
      RECT 671.155 0.155 671.415 13.21 ;
      RECT 669.915 384.61 670.115 385.34 ;
      RECT 670.325 384.61 670.685 385.34 ;
      RECT 670.895 384.61 671.095 385.34 ;
      RECT 671.55 384.61 671.75 385.34 ;
      RECT 671.96 384.61 672.32 385.34 ;
      RECT 672.615 384.61 672.815 385.34 ;
      RECT 673.11 384.61 673.47 385.34 ;
      RECT 673.35 0.52 673.61 14.115 ;
      RECT 673.68 384.61 673.88 385.34 ;
      RECT 673.86 0.52 674.12 13.45 ;
      RECT 674.335 384.61 674.535 385.34 ;
      RECT 674.88 0.155 675.65 0.445 ;
      RECT 674.88 0.155 675.14 8.665 ;
      RECT 675.39 0.155 675.65 8.665 ;
      RECT 674.37 0.52 674.63 11.315 ;
      RECT 674.745 384.61 675.105 385.34 ;
      RECT 675.315 384.61 675.515 385.34 ;
      RECT 675.9 0.52 676.16 9.955 ;
      RECT 675.97 384.61 676.17 385.34 ;
      RECT 676.38 384.61 676.74 385.34 ;
      RECT 677.035 384.61 677.235 385.34 ;
      RECT 677.53 384.61 677.89 385.34 ;
      RECT 677.94 0.3 678.2 8.7 ;
      RECT 678.1 384.61 678.3 385.34 ;
      RECT 678.755 384.61 678.955 385.34 ;
      RECT 678.45 0.18 679.22 0.88 ;
      RECT 679.165 384.61 679.525 385.34 ;
      RECT 679.735 384.61 679.935 385.34 ;
      RECT 680.39 384.61 680.59 385.34 ;
      RECT 680.645 0.52 680.905 6.28 ;
      RECT 680.8 384.61 681.16 385.34 ;
      RECT 681.455 384.61 681.655 385.34 ;
      RECT 682.02 0.52 682.28 5.57 ;
      RECT 681.95 384.61 682.31 385.34 ;
      RECT 682.52 384.61 682.72 385.34 ;
      RECT 682.53 0.3 682.79 5.235 ;
      RECT 683.04 0.52 683.3 7.78 ;
      RECT 683.175 384.61 683.375 385.34 ;
      RECT 683.585 384.61 683.945 385.34 ;
      RECT 684.155 384.61 684.355 385.34 ;
      RECT 684.98 53.41 685.18 385.34 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 681.165 0 681.76 385.37 ;
      RECT 682.53 0.3 682.79 385.37 ;
      RECT 683.56 0 685.49 385.37 ;
      RECT 0 0.52 685.49 385.37 ;
      RECT 676.42 0 680.385 385.37 ;
      RECT 674.88 0.155 675.65 385.37 ;
      RECT 669.435 0 673.09 385.37 ;
      RECT 667.905 0 668.655 385.37 ;
      RECT 666.73 0 667.125 385.37 ;
      RECT 664.85 0.3 665.11 385.37 ;
      RECT 663.485 0 664.08 385.37 ;
      RECT 658.74 0 662.705 385.37 ;
      RECT 657.2 0.155 657.97 385.37 ;
      RECT 651.755 0 655.41 385.37 ;
      RECT 650.225 0 650.975 385.37 ;
      RECT 649.05 0 649.445 385.37 ;
      RECT 647.17 0.3 647.43 385.37 ;
      RECT 645.805 0 646.4 385.37 ;
      RECT 641.06 0 645.025 385.37 ;
      RECT 639.52 0.155 640.29 385.37 ;
      RECT 634.075 0 637.73 385.37 ;
      RECT 632.545 0 633.295 385.37 ;
      RECT 631.37 0 631.765 385.37 ;
      RECT 629.49 0.3 629.75 385.37 ;
      RECT 628.125 0 628.72 385.37 ;
      RECT 623.38 0 627.345 385.37 ;
      RECT 621.84 0.155 622.61 385.37 ;
      RECT 616.395 0 620.05 385.37 ;
      RECT 614.865 0 615.615 385.37 ;
      RECT 613.69 0 614.085 385.37 ;
      RECT 611.81 0.3 612.07 385.37 ;
      RECT 610.445 0 611.04 385.37 ;
      RECT 605.7 0 609.665 385.37 ;
      RECT 604.16 0.155 604.93 385.37 ;
      RECT 598.715 0 602.37 385.37 ;
      RECT 597.185 0 597.935 385.37 ;
      RECT 596.01 0 596.405 385.37 ;
      RECT 594.13 0.3 594.39 385.37 ;
      RECT 592.765 0 593.36 385.37 ;
      RECT 588.02 0 591.985 385.37 ;
      RECT 586.48 0.155 587.25 385.37 ;
      RECT 581.035 0 584.69 385.37 ;
      RECT 579.505 0 580.255 385.37 ;
      RECT 578.33 0 578.725 385.37 ;
      RECT 576.45 0.3 576.71 385.37 ;
      RECT 575.085 0 575.68 385.37 ;
      RECT 570.34 0 574.305 385.37 ;
      RECT 568.8 0.155 569.57 385.37 ;
      RECT 563.355 0 567.01 385.37 ;
      RECT 561.825 0 562.575 385.37 ;
      RECT 560.65 0 561.045 385.37 ;
      RECT 558.77 0.3 559.03 385.37 ;
      RECT 557.405 0 558 385.37 ;
      RECT 552.66 0 556.625 385.37 ;
      RECT 551.12 0.155 551.89 385.37 ;
      RECT 545.675 0 549.33 385.37 ;
      RECT 544.145 0 544.895 385.37 ;
      RECT 542.97 0 543.365 385.37 ;
      RECT 541.09 0.3 541.35 385.37 ;
      RECT 539.725 0 540.32 385.37 ;
      RECT 534.98 0 538.945 385.37 ;
      RECT 533.44 0.155 534.21 385.37 ;
      RECT 527.995 0 531.65 385.37 ;
      RECT 526.465 0 527.215 385.37 ;
      RECT 525.29 0 525.685 385.37 ;
      RECT 523.41 0.3 523.67 385.37 ;
      RECT 522.045 0 522.64 385.37 ;
      RECT 517.3 0 521.265 385.37 ;
      RECT 515.76 0.155 516.53 385.37 ;
      RECT 510.315 0 513.97 385.37 ;
      RECT 508.785 0 509.535 385.37 ;
      RECT 507.61 0 508.005 385.37 ;
      RECT 505.73 0.3 505.99 385.37 ;
      RECT 504.365 0 504.96 385.37 ;
      RECT 499.62 0 503.585 385.37 ;
      RECT 498.08 0.155 498.85 385.37 ;
      RECT 492.635 0 496.29 385.37 ;
      RECT 491.105 0 491.855 385.37 ;
      RECT 489.93 0 490.325 385.37 ;
      RECT 488.05 0.3 488.31 385.37 ;
      RECT 486.685 0 487.28 385.37 ;
      RECT 481.94 0 485.905 385.37 ;
      RECT 480.4 0.155 481.17 385.37 ;
      RECT 474.955 0 478.61 385.37 ;
      RECT 473.425 0 474.175 385.37 ;
      RECT 472.25 0 472.645 385.37 ;
      RECT 470.37 0.3 470.63 385.37 ;
      RECT 469.005 0 469.6 385.37 ;
      RECT 464.26 0 468.225 385.37 ;
      RECT 462.72 0.155 463.49 385.37 ;
      RECT 457.275 0 460.93 385.37 ;
      RECT 455.745 0 456.495 385.37 ;
      RECT 454.57 0 454.965 385.37 ;
      RECT 452.69 0.3 452.95 385.37 ;
      RECT 451.325 0 451.92 385.37 ;
      RECT 446.58 0 450.545 385.37 ;
      RECT 445.04 0.155 445.81 385.37 ;
      RECT 439.595 0 443.25 385.37 ;
      RECT 438.065 0 438.815 385.37 ;
      RECT 436.89 0 437.285 385.37 ;
      RECT 435.01 0.3 435.27 385.37 ;
      RECT 433.645 0 434.24 385.37 ;
      RECT 428.9 0 432.865 385.37 ;
      RECT 427.36 0.155 428.13 385.37 ;
      RECT 421.915 0 425.57 385.37 ;
      RECT 420.385 0 421.135 385.37 ;
      RECT 419.21 0 419.605 385.37 ;
      RECT 417.33 0.3 417.59 385.37 ;
      RECT 415.965 0 416.56 385.37 ;
      RECT 411.22 0 415.185 385.37 ;
      RECT 409.68 0.155 410.45 385.37 ;
      RECT 404.235 0 407.89 385.37 ;
      RECT 402.705 0 403.455 385.37 ;
      RECT 401.53 0 401.925 385.37 ;
      RECT 378.725 0.18 400.75 385.37 ;
      RECT 378.735 0 400.75 385.37 ;
      RECT 374.135 0.3 377.965 385.37 ;
      RECT 372.095 0.18 372.865 385.37 ;
      RECT 365.465 0.3 366.745 385.37 ;
      RECT 362.915 0.3 364.195 385.37 ;
      RECT 361.385 0.3 361.645 385.37 ;
      RECT 358.325 0.3 358.585 385.37 ;
      RECT 356.795 0.3 357.055 385.37 ;
      RECT 348.635 0.3 355.525 385.37 ;
      RECT 339.145 0 346.345 385.37 ;
      RECT 329.965 0.3 336.855 385.37 ;
      RECT 329.975 0 336.855 385.37 ;
      RECT 328.435 0.3 328.695 385.37 ;
      RECT 326.905 0.3 327.165 385.37 ;
      RECT 323.845 0.3 324.105 385.37 ;
      RECT 321.295 0.3 322.575 385.37 ;
      RECT 318.745 0.3 320.025 385.37 ;
      RECT 312.625 0.18 313.395 385.37 ;
      RECT 307.525 0.3 311.355 385.37 ;
      RECT 284.74 0.18 306.765 385.37 ;
      RECT 283.565 0 283.96 385.37 ;
      RECT 282.035 0 282.785 385.37 ;
      RECT 277.6 0 281.255 385.37 ;
      RECT 275.04 0.155 275.81 385.37 ;
      RECT 270.305 0 274.27 385.37 ;
      RECT 268.93 0 269.525 385.37 ;
      RECT 267.9 0.3 268.16 385.37 ;
      RECT 265.885 0 266.28 385.37 ;
      RECT 264.355 0 265.105 385.37 ;
      RECT 259.92 0 263.575 385.37 ;
      RECT 257.36 0.155 258.13 385.37 ;
      RECT 252.625 0 256.59 385.37 ;
      RECT 251.25 0 251.845 385.37 ;
      RECT 250.22 0.3 250.48 385.37 ;
      RECT 248.205 0 248.6 385.37 ;
      RECT 246.675 0 247.425 385.37 ;
      RECT 242.24 0 245.895 385.37 ;
      RECT 239.68 0.155 240.45 385.37 ;
      RECT 234.945 0 238.91 385.37 ;
      RECT 233.57 0 234.165 385.37 ;
      RECT 232.54 0.3 232.8 385.37 ;
      RECT 230.525 0 230.92 385.37 ;
      RECT 228.995 0 229.745 385.37 ;
      RECT 224.56 0 228.215 385.37 ;
      RECT 222 0.155 222.77 385.37 ;
      RECT 217.265 0 221.23 385.37 ;
      RECT 215.89 0 216.485 385.37 ;
      RECT 214.86 0.3 215.12 385.37 ;
      RECT 212.845 0 213.24 385.37 ;
      RECT 211.315 0 212.065 385.37 ;
      RECT 206.88 0 210.535 385.37 ;
      RECT 204.32 0.155 205.09 385.37 ;
      RECT 199.585 0 203.55 385.37 ;
      RECT 198.21 0 198.805 385.37 ;
      RECT 197.18 0.3 197.44 385.37 ;
      RECT 195.165 0 195.56 385.37 ;
      RECT 193.635 0 194.385 385.37 ;
      RECT 189.2 0 192.855 385.37 ;
      RECT 186.64 0.155 187.41 385.37 ;
      RECT 181.905 0 185.87 385.37 ;
      RECT 180.53 0 181.125 385.37 ;
      RECT 179.5 0.3 179.76 385.37 ;
      RECT 177.485 0 177.88 385.37 ;
      RECT 175.955 0 176.705 385.37 ;
      RECT 171.52 0 175.175 385.37 ;
      RECT 168.96 0.155 169.73 385.37 ;
      RECT 164.225 0 168.19 385.37 ;
      RECT 162.85 0 163.445 385.37 ;
      RECT 161.82 0.3 162.08 385.37 ;
      RECT 159.805 0 160.2 385.37 ;
      RECT 158.275 0 159.025 385.37 ;
      RECT 153.84 0 157.495 385.37 ;
      RECT 151.28 0.155 152.05 385.37 ;
      RECT 146.545 0 150.51 385.37 ;
      RECT 145.17 0 145.765 385.37 ;
      RECT 144.14 0.3 144.4 385.37 ;
      RECT 142.125 0 142.52 385.37 ;
      RECT 140.595 0 141.345 385.37 ;
      RECT 136.16 0 139.815 385.37 ;
      RECT 133.6 0.155 134.37 385.37 ;
      RECT 128.865 0 132.83 385.37 ;
      RECT 127.49 0 128.085 385.37 ;
      RECT 126.46 0.3 126.72 385.37 ;
      RECT 124.445 0 124.84 385.37 ;
      RECT 122.915 0 123.665 385.37 ;
      RECT 118.48 0 122.135 385.37 ;
      RECT 115.92 0.155 116.69 385.37 ;
      RECT 111.185 0 115.15 385.37 ;
      RECT 109.81 0 110.405 385.37 ;
      RECT 108.78 0.3 109.04 385.37 ;
      RECT 106.765 0 107.16 385.37 ;
      RECT 105.235 0 105.985 385.37 ;
      RECT 100.8 0 104.455 385.37 ;
      RECT 98.24 0.155 99.01 385.37 ;
      RECT 93.505 0 97.47 385.37 ;
      RECT 92.13 0 92.725 385.37 ;
      RECT 91.1 0.3 91.36 385.37 ;
      RECT 89.085 0 89.48 385.37 ;
      RECT 87.555 0 88.305 385.37 ;
      RECT 83.12 0 86.775 385.37 ;
      RECT 80.56 0.155 81.33 385.37 ;
      RECT 75.825 0 79.79 385.37 ;
      RECT 74.45 0 75.045 385.37 ;
      RECT 73.42 0.3 73.68 385.37 ;
      RECT 71.405 0 71.8 385.37 ;
      RECT 69.875 0 70.625 385.37 ;
      RECT 65.44 0 69.095 385.37 ;
      RECT 62.88 0.155 63.65 385.37 ;
      RECT 58.145 0 62.11 385.37 ;
      RECT 56.77 0 57.365 385.37 ;
      RECT 55.74 0.3 56 385.37 ;
      RECT 53.725 0 54.12 385.37 ;
      RECT 52.195 0 52.945 385.37 ;
      RECT 47.76 0 51.415 385.37 ;
      RECT 45.2 0.155 45.97 385.37 ;
      RECT 40.465 0 44.43 385.37 ;
      RECT 39.09 0 39.685 385.37 ;
      RECT 38.06 0.3 38.32 385.37 ;
      RECT 36.045 0 36.44 385.37 ;
      RECT 34.515 0 35.265 385.37 ;
      RECT 30.08 0 33.735 385.37 ;
      RECT 27.52 0.155 28.29 385.37 ;
      RECT 22.785 0 26.75 385.37 ;
      RECT 21.41 0 22.005 385.37 ;
      RECT 20.38 0.3 20.64 385.37 ;
      RECT 18.365 0 18.76 385.37 ;
      RECT 16.835 0 17.585 385.37 ;
      RECT 12.4 0 16.055 385.37 ;
      RECT 9.84 0.155 10.61 385.37 ;
      RECT 5.105 0 9.07 385.37 ;
      RECT 3.73 0 4.325 385.37 ;
      RECT 2.7 0.3 2.96 385.37 ;
      RECT 0 0 1.93 385.37 ;
      RECT 682.54 0 682.78 385.37 ;
      RECT 664.86 0 665.1 385.37 ;
      RECT 647.18 0 647.42 385.37 ;
      RECT 629.5 0 629.74 385.37 ;
      RECT 611.82 0 612.06 385.37 ;
      RECT 594.14 0 594.38 385.37 ;
      RECT 576.46 0 576.7 385.37 ;
      RECT 558.78 0 559.02 385.37 ;
      RECT 541.1 0 541.34 385.37 ;
      RECT 523.42 0 523.66 385.37 ;
      RECT 505.74 0 505.98 385.37 ;
      RECT 488.06 0 488.3 385.37 ;
      RECT 470.38 0 470.62 385.37 ;
      RECT 452.7 0 452.94 385.37 ;
      RECT 435.02 0 435.26 385.37 ;
      RECT 417.34 0 417.58 385.37 ;
      RECT 374.145 0 377.955 385.37 ;
      RECT 365.475 0 366.735 385.37 ;
      RECT 362.925 0 364.185 385.37 ;
      RECT 361.395 0 361.635 385.37 ;
      RECT 358.335 0 358.575 385.37 ;
      RECT 356.805 0 357.045 385.37 ;
      RECT 348.635 0 355.515 385.37 ;
      RECT 328.445 0 328.685 385.37 ;
      RECT 326.915 0 327.155 385.37 ;
      RECT 323.855 0 324.095 385.37 ;
      RECT 321.305 0 322.565 385.37 ;
      RECT 318.755 0 320.015 385.37 ;
      RECT 307.535 0 311.345 385.37 ;
      RECT 267.91 0 268.15 385.37 ;
      RECT 250.23 0 250.47 385.37 ;
      RECT 232.55 0 232.79 385.37 ;
      RECT 214.87 0 215.11 385.37 ;
      RECT 197.19 0 197.43 385.37 ;
      RECT 179.51 0 179.75 385.37 ;
      RECT 161.83 0 162.07 385.37 ;
      RECT 144.15 0 144.39 385.37 ;
      RECT 126.47 0 126.71 385.37 ;
      RECT 108.79 0 109.03 385.37 ;
      RECT 91.11 0 91.35 385.37 ;
      RECT 73.43 0 73.67 385.37 ;
      RECT 55.75 0 55.99 385.37 ;
      RECT 38.07 0 38.31 385.37 ;
      RECT 20.39 0 20.63 385.37 ;
      RECT 2.71 0 2.95 385.37 ;
      RECT 372.105 0 372.855 385.37 ;
      RECT 312.635 0 313.385 385.37 ;
      RECT 284.74 0 306.755 385.37 ;
      RECT 674.89 0 675.64 385.37 ;
      RECT 657.21 0 657.96 385.37 ;
      RECT 639.53 0 640.28 385.37 ;
      RECT 621.85 0 622.6 385.37 ;
      RECT 604.17 0 604.92 385.37 ;
      RECT 586.49 0 587.24 385.37 ;
      RECT 568.81 0 569.56 385.37 ;
      RECT 551.13 0 551.88 385.37 ;
      RECT 533.45 0 534.2 385.37 ;
      RECT 515.77 0 516.52 385.37 ;
      RECT 498.09 0 498.84 385.37 ;
      RECT 480.41 0 481.16 385.37 ;
      RECT 462.73 0 463.48 385.37 ;
      RECT 445.05 0 445.8 385.37 ;
      RECT 427.37 0 428.12 385.37 ;
      RECT 409.69 0 410.44 385.37 ;
      RECT 275.05 0 275.8 385.37 ;
      RECT 257.37 0 258.12 385.37 ;
      RECT 239.69 0 240.44 385.37 ;
      RECT 222.01 0 222.76 385.37 ;
      RECT 204.33 0 205.08 385.37 ;
      RECT 186.65 0 187.4 385.37 ;
      RECT 168.97 0 169.72 385.37 ;
      RECT 151.29 0 152.04 385.37 ;
      RECT 133.61 0 134.36 385.37 ;
      RECT 115.93 0 116.68 385.37 ;
      RECT 98.25 0 99 385.37 ;
      RECT 80.57 0 81.32 385.37 ;
      RECT 62.89 0 63.64 385.37 ;
      RECT 45.21 0 45.96 385.37 ;
      RECT 27.53 0 28.28 385.37 ;
      RECT 9.85 0 10.6 385.37 ;
    LAYER Metal3 ;
      RECT 0 0 685.49 385.37 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 383.035 0 400.625 385.37 ;
      RECT 377.885 0 379.705 385.37 ;
      RECT 372.735 0 374.555 385.37 ;
      RECT 679.605 0 685.49 385.37 ;
      RECT 670.765 0 674.665 385.37 ;
      RECT 670.765 47.305 685.49 53.15 ;
      RECT 661.925 0 665.825 385.37 ;
      RECT 653.085 0 656.985 385.37 ;
      RECT 653.085 47.305 665.825 53.15 ;
      RECT 644.245 0 648.145 385.37 ;
      RECT 635.405 0 639.305 385.37 ;
      RECT 635.405 47.305 648.145 53.15 ;
      RECT 626.565 0 630.465 385.37 ;
      RECT 617.725 0 621.625 385.37 ;
      RECT 617.725 47.305 630.465 53.15 ;
      RECT 608.885 0 612.785 385.37 ;
      RECT 600.045 0 603.945 385.37 ;
      RECT 600.045 47.305 612.785 53.15 ;
      RECT 591.205 0 595.105 385.37 ;
      RECT 582.365 0 586.265 385.37 ;
      RECT 582.365 47.305 595.105 53.15 ;
      RECT 573.525 0 577.425 385.37 ;
      RECT 564.685 0 568.585 385.37 ;
      RECT 564.685 47.305 577.425 53.15 ;
      RECT 555.845 0 559.745 385.37 ;
      RECT 547.005 0 550.905 385.37 ;
      RECT 547.005 47.305 559.745 53.15 ;
      RECT 538.165 0 542.065 385.37 ;
      RECT 529.325 0 533.225 385.37 ;
      RECT 529.325 47.305 542.065 53.15 ;
      RECT 520.485 0 524.385 385.37 ;
      RECT 511.645 0 515.545 385.37 ;
      RECT 511.645 47.305 524.385 53.15 ;
      RECT 502.805 0 506.705 385.37 ;
      RECT 493.965 0 497.865 385.37 ;
      RECT 493.965 47.305 506.705 53.15 ;
      RECT 485.125 0 489.025 385.37 ;
      RECT 476.285 0 480.185 385.37 ;
      RECT 476.285 47.305 489.025 53.15 ;
      RECT 467.445 0 471.345 385.37 ;
      RECT 458.605 0 462.505 385.37 ;
      RECT 458.605 47.305 471.345 53.15 ;
      RECT 449.765 0 453.665 385.37 ;
      RECT 440.925 0 444.825 385.37 ;
      RECT 440.925 47.305 453.665 53.15 ;
      RECT 432.085 0 435.985 385.37 ;
      RECT 423.245 0 427.145 385.37 ;
      RECT 423.245 47.305 435.985 53.15 ;
      RECT 414.405 0 418.305 385.37 ;
      RECT 405.565 0 409.465 385.37 ;
      RECT 405.565 47.305 418.305 53.15 ;
      RECT 367.585 0 369.405 385.37 ;
      RECT 362.435 0 364.255 385.37 ;
      RECT 357.285 0 359.105 385.37 ;
      RECT 352.135 0 353.955 385.37 ;
      RECT 346.985 0 348.805 385.37 ;
      RECT 341.835 0 343.655 385.37 ;
      RECT 336.685 0 338.505 385.37 ;
      RECT 331.535 0 333.355 385.37 ;
      RECT 326.385 0 328.205 385.37 ;
      RECT 321.235 0 323.055 385.37 ;
      RECT 316.085 0 317.905 385.37 ;
      RECT 310.935 0 312.755 385.37 ;
      RECT 305.785 0 307.605 385.37 ;
      RECT 284.865 0 302.455 385.37 ;
      RECT 276.025 0 279.925 385.37 ;
      RECT 267.185 0 271.085 385.37 ;
      RECT 267.185 47.305 279.925 53.15 ;
      RECT 258.345 0 262.245 385.37 ;
      RECT 249.505 0 253.405 385.37 ;
      RECT 249.505 47.305 262.245 53.15 ;
      RECT 240.665 0 244.565 385.37 ;
      RECT 231.825 0 235.725 385.37 ;
      RECT 231.825 47.305 244.565 53.15 ;
      RECT 222.985 0 226.885 385.37 ;
      RECT 214.145 0 218.045 385.37 ;
      RECT 214.145 47.305 226.885 53.15 ;
      RECT 205.305 0 209.205 385.37 ;
      RECT 196.465 0 200.365 385.37 ;
      RECT 196.465 47.305 209.205 53.15 ;
      RECT 187.625 0 191.525 385.37 ;
      RECT 178.785 0 182.685 385.37 ;
      RECT 178.785 47.305 191.525 53.15 ;
      RECT 169.945 0 173.845 385.37 ;
      RECT 161.105 0 165.005 385.37 ;
      RECT 161.105 47.305 173.845 53.15 ;
      RECT 152.265 0 156.165 385.37 ;
      RECT 143.425 0 147.325 385.37 ;
      RECT 143.425 47.305 156.165 53.15 ;
      RECT 134.585 0 138.485 385.37 ;
      RECT 125.745 0 129.645 385.37 ;
      RECT 125.745 47.305 138.485 53.15 ;
      RECT 116.905 0 120.805 385.37 ;
      RECT 108.065 0 111.965 385.37 ;
      RECT 108.065 47.305 120.805 53.15 ;
      RECT 99.225 0 103.125 385.37 ;
      RECT 90.385 0 94.285 385.37 ;
      RECT 90.385 47.305 103.125 53.15 ;
      RECT 81.545 0 85.445 385.37 ;
      RECT 72.705 0 76.605 385.37 ;
      RECT 72.705 47.305 85.445 53.15 ;
      RECT 63.865 0 67.765 385.37 ;
      RECT 55.025 0 58.925 385.37 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 385.37 ;
      RECT 37.345 0 41.245 385.37 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 385.37 ;
      RECT 19.665 0 23.565 385.37 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 385.37 ;
      RECT 0 0 5.885 385.37 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_1024x32_c2_bm_bist

END LIBRARY
