# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 13:34:44 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_512x8_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_512x8_c2_bm_bist 0 0 ;
  SIZE 261.17 BY 219.77 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.99 0 196.25 0.26 ;
    END
  END A_DIN[4]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.5 0 196.76 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.66 0 204.92 0.26 ;
    END
  END A_BM[4]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.285 0 203.545 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.85 0 189.11 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 198.54 0 198.8 0.26 ;
    END
  END B_DIN[4]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 197.01 0 197.27 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 190.025 0 190.285 0.26 ;
    END
  END B_BM[4]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 191.555 0 191.815 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.68 0 205.94 0.26 ;
    END
  END B_DOUT[4]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 241.765 0 246.185 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.085 0 228.505 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.405 0 210.825 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 188.725 0 193.145 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.805 0 170.615 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 157.505 0 160.315 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 142.055 0 144.865 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 131.755 0 134.565 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.605 0 129.415 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.305 0 119.115 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 100.855 0 103.665 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.555 0 93.365 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 219.77 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 250.605 0 255.025 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 232.925 0 237.345 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.245 0 219.665 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 197.565 0 201.985 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.655 0 165.465 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 152.355 0 155.165 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.205 0 150.015 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 136.905 0 139.715 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.455 0 124.265 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.155 0 113.965 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.005 0 108.815 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 95.705 0 98.515 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 250.605 53.41 255.025 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 232.925 53.41 237.345 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 215.245 53.41 219.665 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 197.565 53.41 201.985 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 219.77 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 219.77 ;
    END
  END VDDARRAY!
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.67 0 213.93 0.26 ;
    END
  END A_DIN[5]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.18 0 214.44 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 222.34 0 222.6 0.26 ;
    END
  END A_BM[5]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 220.965 0 221.225 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.53 0 206.79 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 216.22 0 216.48 0.26 ;
    END
  END B_DIN[5]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.69 0 214.95 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.705 0 207.965 0.26 ;
    END
  END B_BM[5]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 209.235 0 209.495 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.36 0 223.62 0.26 ;
    END
  END B_DOUT[5]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.35 0 231.61 0.26 ;
    END
  END A_DIN[6]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.86 0 232.12 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 240.02 0 240.28 0.26 ;
    END
  END A_BM[6]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 238.645 0 238.905 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.21 0 224.47 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 233.9 0 234.16 0.26 ;
    END
  END B_DIN[6]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.37 0 232.63 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 225.385 0 225.645 0.26 ;
    END
  END B_BM[6]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.915 0 227.175 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.04 0 241.3 0.26 ;
    END
  END B_DOUT[6]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.03 0 249.29 0.26 ;
    END
  END A_DIN[7]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.54 0 249.8 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 257.7 0 257.96 0.26 ;
    END
  END A_BM[7]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 256.325 0 256.585 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.89 0 242.15 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 251.58 0 251.84 0.26 ;
    END
  END B_DIN[7]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 250.05 0 250.31 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 243.065 0 243.325 0.26 ;
    END
  END B_BM[7]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 244.595 0 244.855 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.72 0 258.98 0.26 ;
    END
  END B_DOUT[7]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.675 0 146.935 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.285 0 152.545 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.235 0 114.495 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.625 0 108.885 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 147.185 0 147.445 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.795 0 153.055 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.725 0 113.985 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.115 0 108.375 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 155.855 0 156.115 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 156.365 0 156.625 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 105.055 0 105.315 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 104.545 0 104.805 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 154.835 0 155.095 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 155.345 0 155.605 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 106.075 0 106.335 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 105.565 0 105.825 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.455 0 135.715 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.965 0 136.225 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.455 0 125.715 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.945 0 125.205 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.435 0 134.695 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.945 0 135.205 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.475 0 126.735 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.965 0 126.225 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.405 0 158.665 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.895 0 158.155 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.505 0 102.765 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.015 0 103.275 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.385 0 157.645 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.875 0 157.135 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.525 0 103.785 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.035 0 104.295 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.955 0 161.215 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.465 0 161.725 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN B_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4422 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.811551 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.955 0 100.215 0.26 ;
    END
  END B_ADDR[8]
  PIN B_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.541947 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.445 0 99.705 0.26 ;
    END
  END B_BIST_ADDR[8]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.145 0 145.405 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 148.715 0 148.975 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 148.205 0 148.465 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.655 0 145.915 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 166.055 0 166.315 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.765 0 116.025 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.195 0 112.455 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.705 0 112.965 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.255 0 115.515 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 94.855 0 95.115 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 92.8757 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.3675 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.129726 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 147.695 0 147.955 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.615 0 143.875 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.245 0 150.505 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 149.735 0 149.995 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.125 0 144.385 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 93.3149 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.3675 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.172089 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.215 0 113.475 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.295 0 117.555 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.665 0 110.925 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.175 0 111.435 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.785 0 117.045 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 261.17 219.77 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 219.74 ;
      RECT 1.135 219.01 1.335 219.74 ;
      RECT 1.545 219.01 1.905 219.74 ;
      RECT 2.115 219.01 2.315 219.74 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 219.01 2.97 219.74 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 219.01 3.54 219.74 ;
      RECT 3.835 219.01 4.035 219.74 ;
      RECT 4.33 219.01 4.69 219.74 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 219.01 5.1 219.74 ;
      RECT 5.555 219.01 5.755 219.74 ;
      RECT 5.965 219.01 6.325 219.74 ;
      RECT 6.535 219.01 6.735 219.74 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 219.01 7.39 219.74 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 219.01 7.96 219.74 ;
      RECT 8.255 219.01 8.455 219.74 ;
      RECT 8.75 219.01 9.11 219.74 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 219.01 9.52 219.74 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 219.01 10.175 219.74 ;
      RECT 10.385 219.01 10.745 219.74 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 219.01 11.155 219.74 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 219.01 11.81 219.74 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 219.01 12.38 219.74 ;
      RECT 12.675 219.01 12.875 219.74 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 219.01 13.53 219.74 ;
      RECT 13.74 219.01 13.94 219.74 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 219.01 14.595 219.74 ;
      RECT 14.805 219.01 15.165 219.74 ;
      RECT 15.375 219.01 15.575 219.74 ;
      RECT 16.03 219.01 16.23 219.74 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 219.01 16.8 219.74 ;
      RECT 17.095 219.01 17.295 219.74 ;
      RECT 17.59 219.01 17.95 219.74 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 219.01 18.36 219.74 ;
      RECT 18.815 219.01 19.015 219.74 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 219.01 19.585 219.74 ;
      RECT 19.795 219.01 19.995 219.74 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 219.01 20.65 219.74 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 219.01 21.22 219.74 ;
      RECT 21.515 219.01 21.715 219.74 ;
      RECT 22.01 219.01 22.37 219.74 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 219.01 22.78 219.74 ;
      RECT 23.235 219.01 23.435 219.74 ;
      RECT 23.645 219.01 24.005 219.74 ;
      RECT 24.215 219.01 24.415 219.74 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 219.01 25.07 219.74 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 219.01 25.64 219.74 ;
      RECT 25.935 219.01 26.135 219.74 ;
      RECT 26.43 219.01 26.79 219.74 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 219.01 27.2 219.74 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 219.01 27.855 219.74 ;
      RECT 28.065 219.01 28.425 219.74 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 219.01 28.835 219.74 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 219.01 29.49 219.74 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 219.01 30.06 219.74 ;
      RECT 30.355 219.01 30.555 219.74 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 219.01 31.21 219.74 ;
      RECT 31.42 219.01 31.62 219.74 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 219.01 32.275 219.74 ;
      RECT 32.485 219.01 32.845 219.74 ;
      RECT 33.055 219.01 33.255 219.74 ;
      RECT 33.71 219.01 33.91 219.74 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 219.01 34.48 219.74 ;
      RECT 34.775 219.01 34.975 219.74 ;
      RECT 35.27 219.01 35.63 219.74 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 219.01 36.04 219.74 ;
      RECT 36.495 219.01 36.695 219.74 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 219.01 37.265 219.74 ;
      RECT 37.475 219.01 37.675 219.74 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 219.01 38.33 219.74 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 219.01 38.9 219.74 ;
      RECT 39.195 219.01 39.395 219.74 ;
      RECT 39.69 219.01 40.05 219.74 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 219.01 40.46 219.74 ;
      RECT 40.915 219.01 41.115 219.74 ;
      RECT 41.325 219.01 41.685 219.74 ;
      RECT 41.895 219.01 42.095 219.74 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 219.01 42.75 219.74 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 219.01 43.32 219.74 ;
      RECT 43.615 219.01 43.815 219.74 ;
      RECT 44.11 219.01 44.47 219.74 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 219.01 44.88 219.74 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 219.01 45.535 219.74 ;
      RECT 45.745 219.01 46.105 219.74 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 219.01 46.515 219.74 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 219.01 47.17 219.74 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 219.01 47.74 219.74 ;
      RECT 48.035 219.01 48.235 219.74 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 219.01 48.89 219.74 ;
      RECT 49.1 219.01 49.3 219.74 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 219.01 49.955 219.74 ;
      RECT 50.165 219.01 50.525 219.74 ;
      RECT 50.735 219.01 50.935 219.74 ;
      RECT 51.39 219.01 51.59 219.74 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 219.01 52.16 219.74 ;
      RECT 52.455 219.01 52.655 219.74 ;
      RECT 52.95 219.01 53.31 219.74 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 219.01 53.72 219.74 ;
      RECT 54.175 219.01 54.375 219.74 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 219.01 54.945 219.74 ;
      RECT 55.155 219.01 55.355 219.74 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 219.01 56.01 219.74 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 219.01 56.58 219.74 ;
      RECT 56.875 219.01 57.075 219.74 ;
      RECT 57.37 219.01 57.73 219.74 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 219.01 58.14 219.74 ;
      RECT 58.595 219.01 58.795 219.74 ;
      RECT 59.005 219.01 59.365 219.74 ;
      RECT 59.575 219.01 59.775 219.74 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 219.01 60.43 219.74 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 219.01 61 219.74 ;
      RECT 61.295 219.01 61.495 219.74 ;
      RECT 61.79 219.01 62.15 219.74 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 219.01 62.56 219.74 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 219.01 63.215 219.74 ;
      RECT 63.425 219.01 63.785 219.74 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 219.01 64.195 219.74 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 219.01 64.85 219.74 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 219.01 65.42 219.74 ;
      RECT 65.715 219.01 65.915 219.74 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 219.01 66.57 219.74 ;
      RECT 66.78 219.01 66.98 219.74 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 219.01 67.635 219.74 ;
      RECT 67.845 219.01 68.205 219.74 ;
      RECT 68.415 219.01 68.615 219.74 ;
      RECT 69.07 219.01 69.27 219.74 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 219.01 69.84 219.74 ;
      RECT 70.135 219.01 70.335 219.74 ;
      RECT 70.63 219.01 70.99 219.74 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 219.01 71.4 219.74 ;
      RECT 71.855 219.01 72.055 219.74 ;
      RECT 73.08 0.17 73.85 0.43 ;
      RECT 73.08 0.17 73.34 8.7 ;
      RECT 73.59 0.17 73.85 8.7 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 74.1 0.18 74.87 0.88 ;
      RECT 74.1 0.18 74.36 8.7 ;
      RECT 74.61 0.18 74.87 8.7 ;
      RECT 75.12 0.17 75.89 0.43 ;
      RECT 75.12 0.17 75.38 8.7 ;
      RECT 75.63 0.17 75.89 8.7 ;
      RECT 76.14 0.18 76.91 0.88 ;
      RECT 76.14 0.18 76.4 8.7 ;
      RECT 76.65 0.18 76.91 8.7 ;
      RECT 77.16 0.17 77.93 0.43 ;
      RECT 77.16 0.17 77.42 8.7 ;
      RECT 77.67 0.17 77.93 8.7 ;
      RECT 78.18 0.18 78.95 0.88 ;
      RECT 78.18 0.18 78.44 8.7 ;
      RECT 78.69 0.18 78.95 8.7 ;
      RECT 79.2 0.17 79.97 0.43 ;
      RECT 79.2 0.17 79.46 8.7 ;
      RECT 79.71 0.17 79.97 8.7 ;
      RECT 80.22 0.18 80.99 0.88 ;
      RECT 80.22 0.18 80.48 8.7 ;
      RECT 80.73 0.18 80.99 8.7 ;
      RECT 81.24 0.17 82.01 0.43 ;
      RECT 81.24 0.17 81.5 8.7 ;
      RECT 81.75 0.17 82.01 8.7 ;
      RECT 82.26 0.18 83.03 0.88 ;
      RECT 82.26 0.18 82.52 8.7 ;
      RECT 82.77 0.18 83.03 8.7 ;
      RECT 83.28 0.17 84.05 0.43 ;
      RECT 83.28 0.17 83.54 8.7 ;
      RECT 83.79 0.17 84.05 8.7 ;
      RECT 84.3 0.18 85.07 0.88 ;
      RECT 84.3 0.18 84.56 8.7 ;
      RECT 84.81 0.18 85.07 8.7 ;
      RECT 85.32 0.17 86.09 0.43 ;
      RECT 85.32 0.17 85.58 8.7 ;
      RECT 85.83 0.17 86.09 8.7 ;
      RECT 86.34 0.18 87.11 0.88 ;
      RECT 86.34 0.18 86.6 8.7 ;
      RECT 86.85 0.18 87.11 8.7 ;
      RECT 87.36 0.17 88.13 0.43 ;
      RECT 87.36 0.17 87.62 8.7 ;
      RECT 87.87 0.17 88.13 8.7 ;
      RECT 88.38 0.18 89.15 0.88 ;
      RECT 88.38 0.18 88.64 8.7 ;
      RECT 88.89 0.18 89.15 8.7 ;
      RECT 72.265 219.01 72.625 219.74 ;
      RECT 72.835 219.01 73.035 219.74 ;
      RECT 90.775 0.18 91.545 0.88 ;
      RECT 90.775 0.18 91.035 8.7 ;
      RECT 91.285 0.18 91.545 8.7 ;
      RECT 91.795 0.17 92.565 0.43 ;
      RECT 91.795 0.17 92.055 8.7 ;
      RECT 92.305 0.17 92.565 8.7 ;
      RECT 73.66 218.93 73.86 219.74 ;
      RECT 89.755 0.3 90.015 8.7 ;
      RECT 93.835 0.18 94.605 0.88 ;
      RECT 93.835 0.18 94.095 8.7 ;
      RECT 94.345 0.18 94.605 8.7 ;
      RECT 90.265 0.3 90.525 8.7 ;
      RECT 92.815 0 93.075 8.7 ;
      RECT 93.325 0 93.585 8.7 ;
      RECT 94.855 0.52 95.115 8.7 ;
      RECT 95.365 0.3 95.625 8.7 ;
      RECT 95.875 0.3 96.135 8.7 ;
      RECT 96.385 0.3 96.645 8.7 ;
      RECT 96.895 0.3 97.155 8.7 ;
      RECT 97.405 0.3 97.665 8.7 ;
      RECT 97.915 0.3 98.175 8.7 ;
      RECT 98.425 0.3 98.685 8.7 ;
      RECT 100.465 0.18 101.235 0.88 ;
      RECT 100.465 0.18 100.725 8.7 ;
      RECT 100.975 0.18 101.235 8.7 ;
      RECT 98.935 0.3 99.195 8.7 ;
      RECT 99.445 0.52 99.705 8.7 ;
      RECT 99.955 0.52 100.215 8.7 ;
      RECT 101.485 0 101.745 8.7 ;
      RECT 101.995 0 102.255 8.7 ;
      RECT 102.505 0.52 102.765 8.7 ;
      RECT 103.015 0.52 103.275 8.7 ;
      RECT 103.525 0.52 103.785 8.7 ;
      RECT 104.035 0.52 104.295 8.7 ;
      RECT 104.545 0.52 104.805 8.7 ;
      RECT 105.055 0.52 105.315 8.7 ;
      RECT 105.565 0.52 105.825 8.7 ;
      RECT 106.075 0.52 106.335 8.7 ;
      RECT 106.585 0.3 106.845 8.7 ;
      RECT 107.095 0.3 107.355 8.7 ;
      RECT 107.605 0.3 107.865 8.7 ;
      RECT 108.115 0.52 108.375 8.7 ;
      RECT 108.625 0.52 108.885 8.7 ;
      RECT 109.135 0.3 109.395 8.7 ;
      RECT 109.645 0.3 109.905 8.7 ;
      RECT 110.155 0.3 110.415 8.7 ;
      RECT 110.665 0.52 110.925 8.7 ;
      RECT 111.175 0.52 111.435 8.7 ;
      RECT 111.685 0.3 111.945 8.7 ;
      RECT 112.195 0.52 112.455 8.7 ;
      RECT 112.705 0.52 112.965 8.7 ;
      RECT 113.215 0.52 113.475 8.7 ;
      RECT 113.725 0.52 113.985 8.7 ;
      RECT 114.235 0.52 114.495 8.7 ;
      RECT 114.745 0.3 115.005 8.7 ;
      RECT 115.255 0.52 115.515 8.7 ;
      RECT 115.765 0.52 116.025 8.7 ;
      RECT 116.275 0.3 116.535 8.7 ;
      RECT 116.785 0.52 117.045 8.7 ;
      RECT 118.825 0.17 119.595 0.43 ;
      RECT 118.825 0.17 119.085 8.7 ;
      RECT 119.335 0.17 119.595 8.7 ;
      RECT 117.295 0.52 117.555 8.7 ;
      RECT 117.805 0.3 118.065 8.7 ;
      RECT 118.315 0.3 118.575 8.7 ;
      RECT 121.375 0.17 122.145 0.43 ;
      RECT 121.375 0.17 121.635 8.7 ;
      RECT 121.885 0.17 122.145 8.7 ;
      RECT 119.845 0.3 120.105 8.7 ;
      RECT 122.905 0.18 123.675 0.88 ;
      RECT 122.905 0.18 123.165 8.7 ;
      RECT 123.415 0.18 123.675 8.7 ;
      RECT 120.355 0.3 120.615 8.7 ;
      RECT 120.865 0.3 121.125 8.7 ;
      RECT 122.395 0.3 122.655 8.7 ;
      RECT 123.925 0 124.185 8.7 ;
      RECT 124.435 0 124.695 8.7 ;
      RECT 124.945 0.52 125.205 8.7 ;
      RECT 125.455 0.52 125.715 8.7 ;
      RECT 125.965 0.52 126.225 8.7 ;
      RECT 126.475 0.52 126.735 8.7 ;
      RECT 126.985 0 127.245 8.7 ;
      RECT 127.495 0 127.755 8.7 ;
      RECT 128.005 0.3 128.265 8.7 ;
      RECT 128.515 0.3 128.775 8.7 ;
      RECT 129.025 0 129.285 8.7 ;
      RECT 129.535 0 129.795 8.7 ;
      RECT 130.045 0.3 130.305 8.7 ;
      RECT 130.865 0.3 131.125 8.7 ;
      RECT 131.375 0 131.635 8.7 ;
      RECT 131.885 0 132.145 8.7 ;
      RECT 132.395 0.3 132.655 8.7 ;
      RECT 132.905 0.3 133.165 8.7 ;
      RECT 133.415 0 133.675 8.7 ;
      RECT 133.925 0 134.185 8.7 ;
      RECT 134.435 0.52 134.695 8.7 ;
      RECT 134.945 0.52 135.205 8.7 ;
      RECT 135.455 0.52 135.715 8.7 ;
      RECT 137.495 0.18 138.265 0.88 ;
      RECT 137.495 0.18 137.755 8.7 ;
      RECT 138.005 0.18 138.265 8.7 ;
      RECT 135.965 0.52 136.225 8.7 ;
      RECT 139.025 0.17 139.795 0.43 ;
      RECT 139.025 0.17 139.285 8.7 ;
      RECT 139.535 0.17 139.795 8.7 ;
      RECT 136.475 0 136.735 8.7 ;
      RECT 136.985 0 137.245 8.7 ;
      RECT 138.515 0.3 138.775 8.7 ;
      RECT 141.575 0.17 142.345 0.43 ;
      RECT 141.575 0.17 141.835 8.7 ;
      RECT 142.085 0.17 142.345 8.7 ;
      RECT 140.045 0.3 140.305 8.7 ;
      RECT 140.555 0.3 140.815 8.7 ;
      RECT 141.065 0.3 141.325 8.7 ;
      RECT 142.595 0.3 142.855 8.7 ;
      RECT 143.105 0.3 143.365 8.7 ;
      RECT 143.615 0.52 143.875 8.7 ;
      RECT 144.125 0.52 144.385 8.7 ;
      RECT 144.635 0.3 144.895 8.7 ;
      RECT 145.145 0.52 145.405 8.7 ;
      RECT 145.655 0.52 145.915 8.7 ;
      RECT 146.165 0.3 146.425 8.7 ;
      RECT 146.675 0.52 146.935 8.7 ;
      RECT 147.185 0.52 147.445 8.7 ;
      RECT 147.695 0.52 147.955 8.7 ;
      RECT 148.205 0.52 148.465 8.7 ;
      RECT 148.715 0.52 148.975 8.7 ;
      RECT 149.225 0.3 149.485 8.7 ;
      RECT 149.735 0.52 149.995 8.7 ;
      RECT 150.245 0.52 150.505 8.7 ;
      RECT 150.755 0.3 151.015 8.7 ;
      RECT 151.265 0.3 151.525 8.7 ;
      RECT 151.775 0.3 152.035 8.7 ;
      RECT 152.285 0.52 152.545 8.7 ;
      RECT 152.795 0.52 153.055 8.7 ;
      RECT 153.305 0.3 153.565 8.7 ;
      RECT 153.815 0.3 154.075 8.7 ;
      RECT 154.325 0.3 154.585 8.7 ;
      RECT 154.835 0.52 155.095 8.7 ;
      RECT 155.345 0.52 155.605 8.7 ;
      RECT 155.855 0.52 156.115 8.7 ;
      RECT 156.365 0.52 156.625 8.7 ;
      RECT 156.875 0.52 157.135 8.7 ;
      RECT 157.385 0.52 157.645 8.7 ;
      RECT 157.895 0.52 158.155 8.7 ;
      RECT 159.935 0.18 160.705 0.88 ;
      RECT 159.935 0.18 160.195 8.7 ;
      RECT 160.445 0.18 160.705 8.7 ;
      RECT 158.405 0.52 158.665 8.7 ;
      RECT 158.915 0 159.175 8.7 ;
      RECT 159.425 0 159.685 8.7 ;
      RECT 160.955 0.52 161.215 8.7 ;
      RECT 161.465 0.52 161.725 8.7 ;
      RECT 161.975 0.3 162.235 8.7 ;
      RECT 162.485 0.3 162.745 8.7 ;
      RECT 162.995 0.3 163.255 8.7 ;
      RECT 163.505 0.3 163.765 8.7 ;
      RECT 164.015 0.3 164.275 8.7 ;
      RECT 164.525 0.3 164.785 8.7 ;
      RECT 166.565 0.18 167.335 0.88 ;
      RECT 166.565 0.18 166.825 8.7 ;
      RECT 167.075 0.18 167.335 8.7 ;
      RECT 165.035 0.3 165.295 8.7 ;
      RECT 165.545 0.3 165.805 8.7 ;
      RECT 168.605 0.17 169.375 0.43 ;
      RECT 168.605 0.17 168.865 8.7 ;
      RECT 169.115 0.17 169.375 8.7 ;
      RECT 169.625 0.18 170.395 0.88 ;
      RECT 169.625 0.18 169.885 8.7 ;
      RECT 170.135 0.18 170.395 8.7 ;
      RECT 166.055 0.52 166.315 8.7 ;
      RECT 167.585 0 167.845 8.7 ;
      RECT 172.02 0.18 172.79 0.88 ;
      RECT 172.02 0.18 172.28 8.7 ;
      RECT 172.53 0.18 172.79 8.7 ;
      RECT 173.04 0.17 173.81 0.43 ;
      RECT 173.04 0.17 173.3 8.7 ;
      RECT 173.55 0.17 173.81 8.7 ;
      RECT 174.06 0.18 174.83 0.88 ;
      RECT 174.06 0.18 174.32 8.7 ;
      RECT 174.57 0.18 174.83 8.7 ;
      RECT 175.08 0.17 175.85 0.43 ;
      RECT 175.08 0.17 175.34 8.7 ;
      RECT 175.59 0.17 175.85 8.7 ;
      RECT 176.1 0.18 176.87 0.88 ;
      RECT 176.1 0.18 176.36 8.7 ;
      RECT 176.61 0.18 176.87 8.7 ;
      RECT 177.12 0.17 177.89 0.43 ;
      RECT 177.12 0.17 177.38 8.7 ;
      RECT 177.63 0.17 177.89 8.7 ;
      RECT 178.14 0.18 178.91 0.88 ;
      RECT 178.14 0.18 178.4 8.7 ;
      RECT 178.65 0.18 178.91 8.7 ;
      RECT 179.16 0.17 179.93 0.43 ;
      RECT 179.16 0.17 179.42 8.7 ;
      RECT 179.67 0.17 179.93 8.7 ;
      RECT 180.18 0.18 180.95 0.88 ;
      RECT 180.18 0.18 180.44 8.7 ;
      RECT 180.69 0.18 180.95 8.7 ;
      RECT 181.2 0.17 181.97 0.43 ;
      RECT 181.2 0.17 181.46 8.7 ;
      RECT 181.71 0.17 181.97 8.7 ;
      RECT 182.22 0.18 182.99 0.88 ;
      RECT 182.22 0.18 182.48 8.7 ;
      RECT 182.73 0.18 182.99 8.7 ;
      RECT 183.24 0.17 184.01 0.43 ;
      RECT 183.24 0.17 183.5 8.7 ;
      RECT 183.75 0.17 184.01 8.7 ;
      RECT 184.26 0.18 185.03 0.88 ;
      RECT 184.26 0.18 184.52 8.7 ;
      RECT 184.77 0.18 185.03 8.7 ;
      RECT 185.28 0.17 186.05 0.43 ;
      RECT 185.28 0.17 185.54 8.7 ;
      RECT 185.79 0.17 186.05 8.7 ;
      RECT 186.3 0.18 187.07 0.88 ;
      RECT 186.3 0.18 186.56 8.7 ;
      RECT 186.81 0.18 187.07 8.7 ;
      RECT 168.095 0 168.355 8.7 ;
      RECT 187.32 0.17 188.09 0.43 ;
      RECT 187.32 0.17 187.58 8.7 ;
      RECT 187.83 0.17 188.09 8.7 ;
      RECT 170.645 0.3 170.905 8.7 ;
      RECT 171.155 0.3 171.415 8.7 ;
      RECT 187.31 218.93 187.51 219.74 ;
      RECT 188.135 219.01 188.335 219.74 ;
      RECT 188.545 219.01 188.905 219.74 ;
      RECT 188.85 0.52 189.11 4.315 ;
      RECT 189.115 219.01 189.315 219.74 ;
      RECT 189.77 219.01 189.97 219.74 ;
      RECT 190.025 0.52 190.285 2.82 ;
      RECT 190.18 219.01 190.54 219.74 ;
      RECT 190.835 219.01 191.035 219.74 ;
      RECT 191.33 219.01 191.69 219.74 ;
      RECT 192.265 0.18 193.035 0.88 ;
      RECT 192.265 0.18 192.525 12.9 ;
      RECT 192.775 0.18 193.035 12.9 ;
      RECT 191.555 0.52 191.815 2.82 ;
      RECT 191.9 219.01 192.1 219.74 ;
      RECT 193.285 0.155 194.055 0.445 ;
      RECT 193.285 0.155 193.545 13.21 ;
      RECT 193.795 0.155 194.055 13.21 ;
      RECT 192.555 219.01 192.755 219.74 ;
      RECT 192.965 219.01 193.325 219.74 ;
      RECT 193.535 219.01 193.735 219.74 ;
      RECT 194.19 219.01 194.39 219.74 ;
      RECT 194.6 219.01 194.96 219.74 ;
      RECT 195.255 219.01 195.455 219.74 ;
      RECT 195.75 219.01 196.11 219.74 ;
      RECT 195.99 0.52 196.25 14.115 ;
      RECT 196.32 219.01 196.52 219.74 ;
      RECT 196.5 0.52 196.76 13.45 ;
      RECT 196.975 219.01 197.175 219.74 ;
      RECT 197.52 0.155 198.29 0.445 ;
      RECT 197.52 0.155 197.78 8.665 ;
      RECT 198.03 0.155 198.29 8.665 ;
      RECT 197.01 0.52 197.27 11.315 ;
      RECT 197.385 219.01 197.745 219.74 ;
      RECT 197.955 219.01 198.155 219.74 ;
      RECT 198.54 0.52 198.8 9.955 ;
      RECT 198.61 219.01 198.81 219.74 ;
      RECT 199.02 219.01 199.38 219.74 ;
      RECT 199.675 219.01 199.875 219.74 ;
      RECT 200.17 219.01 200.53 219.74 ;
      RECT 200.58 0.3 200.84 8.7 ;
      RECT 200.74 219.01 200.94 219.74 ;
      RECT 201.395 219.01 201.595 219.74 ;
      RECT 201.09 0.18 201.86 0.88 ;
      RECT 201.805 219.01 202.165 219.74 ;
      RECT 202.375 219.01 202.575 219.74 ;
      RECT 203.03 219.01 203.23 219.74 ;
      RECT 203.285 0.52 203.545 6.28 ;
      RECT 203.44 219.01 203.8 219.74 ;
      RECT 204.095 219.01 204.295 219.74 ;
      RECT 204.66 0.52 204.92 5.57 ;
      RECT 204.59 219.01 204.95 219.74 ;
      RECT 205.16 219.01 205.36 219.74 ;
      RECT 205.17 0.3 205.43 5.235 ;
      RECT 205.68 0.52 205.94 7.78 ;
      RECT 205.815 219.01 206.015 219.74 ;
      RECT 206.225 219.01 206.585 219.74 ;
      RECT 206.53 0.52 206.79 4.315 ;
      RECT 206.795 219.01 206.995 219.74 ;
      RECT 207.45 219.01 207.65 219.74 ;
      RECT 207.705 0.52 207.965 2.82 ;
      RECT 207.86 219.01 208.22 219.74 ;
      RECT 208.515 219.01 208.715 219.74 ;
      RECT 209.01 219.01 209.37 219.74 ;
      RECT 209.945 0.18 210.715 0.88 ;
      RECT 209.945 0.18 210.205 12.9 ;
      RECT 210.455 0.18 210.715 12.9 ;
      RECT 209.235 0.52 209.495 2.82 ;
      RECT 209.58 219.01 209.78 219.74 ;
      RECT 210.965 0.155 211.735 0.445 ;
      RECT 210.965 0.155 211.225 13.21 ;
      RECT 211.475 0.155 211.735 13.21 ;
      RECT 210.235 219.01 210.435 219.74 ;
      RECT 210.645 219.01 211.005 219.74 ;
      RECT 211.215 219.01 211.415 219.74 ;
      RECT 211.87 219.01 212.07 219.74 ;
      RECT 212.28 219.01 212.64 219.74 ;
      RECT 212.935 219.01 213.135 219.74 ;
      RECT 213.43 219.01 213.79 219.74 ;
      RECT 213.67 0.52 213.93 14.115 ;
      RECT 214 219.01 214.2 219.74 ;
      RECT 214.18 0.52 214.44 13.45 ;
      RECT 214.655 219.01 214.855 219.74 ;
      RECT 215.2 0.155 215.97 0.445 ;
      RECT 215.2 0.155 215.46 8.665 ;
      RECT 215.71 0.155 215.97 8.665 ;
      RECT 214.69 0.52 214.95 11.315 ;
      RECT 215.065 219.01 215.425 219.74 ;
      RECT 215.635 219.01 215.835 219.74 ;
      RECT 216.22 0.52 216.48 9.955 ;
      RECT 216.29 219.01 216.49 219.74 ;
      RECT 216.7 219.01 217.06 219.74 ;
      RECT 217.355 219.01 217.555 219.74 ;
      RECT 217.85 219.01 218.21 219.74 ;
      RECT 218.26 0.3 218.52 8.7 ;
      RECT 218.42 219.01 218.62 219.74 ;
      RECT 219.075 219.01 219.275 219.74 ;
      RECT 218.77 0.18 219.54 0.88 ;
      RECT 219.485 219.01 219.845 219.74 ;
      RECT 220.055 219.01 220.255 219.74 ;
      RECT 220.71 219.01 220.91 219.74 ;
      RECT 220.965 0.52 221.225 6.28 ;
      RECT 221.12 219.01 221.48 219.74 ;
      RECT 221.775 219.01 221.975 219.74 ;
      RECT 222.34 0.52 222.6 5.57 ;
      RECT 222.27 219.01 222.63 219.74 ;
      RECT 222.84 219.01 223.04 219.74 ;
      RECT 222.85 0.3 223.11 5.235 ;
      RECT 223.36 0.52 223.62 7.78 ;
      RECT 223.495 219.01 223.695 219.74 ;
      RECT 223.905 219.01 224.265 219.74 ;
      RECT 224.21 0.52 224.47 4.315 ;
      RECT 224.475 219.01 224.675 219.74 ;
      RECT 225.13 219.01 225.33 219.74 ;
      RECT 225.385 0.52 225.645 2.82 ;
      RECT 225.54 219.01 225.9 219.74 ;
      RECT 226.195 219.01 226.395 219.74 ;
      RECT 226.69 219.01 227.05 219.74 ;
      RECT 227.625 0.18 228.395 0.88 ;
      RECT 227.625 0.18 227.885 12.9 ;
      RECT 228.135 0.18 228.395 12.9 ;
      RECT 226.915 0.52 227.175 2.82 ;
      RECT 227.26 219.01 227.46 219.74 ;
      RECT 228.645 0.155 229.415 0.445 ;
      RECT 228.645 0.155 228.905 13.21 ;
      RECT 229.155 0.155 229.415 13.21 ;
      RECT 227.915 219.01 228.115 219.74 ;
      RECT 228.325 219.01 228.685 219.74 ;
      RECT 228.895 219.01 229.095 219.74 ;
      RECT 229.55 219.01 229.75 219.74 ;
      RECT 229.96 219.01 230.32 219.74 ;
      RECT 230.615 219.01 230.815 219.74 ;
      RECT 231.11 219.01 231.47 219.74 ;
      RECT 231.35 0.52 231.61 14.115 ;
      RECT 231.68 219.01 231.88 219.74 ;
      RECT 231.86 0.52 232.12 13.45 ;
      RECT 232.335 219.01 232.535 219.74 ;
      RECT 232.88 0.155 233.65 0.445 ;
      RECT 232.88 0.155 233.14 8.665 ;
      RECT 233.39 0.155 233.65 8.665 ;
      RECT 232.37 0.52 232.63 11.315 ;
      RECT 232.745 219.01 233.105 219.74 ;
      RECT 233.315 219.01 233.515 219.74 ;
      RECT 233.9 0.52 234.16 9.955 ;
      RECT 233.97 219.01 234.17 219.74 ;
      RECT 234.38 219.01 234.74 219.74 ;
      RECT 235.035 219.01 235.235 219.74 ;
      RECT 235.53 219.01 235.89 219.74 ;
      RECT 235.94 0.3 236.2 8.7 ;
      RECT 236.1 219.01 236.3 219.74 ;
      RECT 236.755 219.01 236.955 219.74 ;
      RECT 236.45 0.18 237.22 0.88 ;
      RECT 237.165 219.01 237.525 219.74 ;
      RECT 237.735 219.01 237.935 219.74 ;
      RECT 238.39 219.01 238.59 219.74 ;
      RECT 238.645 0.52 238.905 6.28 ;
      RECT 238.8 219.01 239.16 219.74 ;
      RECT 239.455 219.01 239.655 219.74 ;
      RECT 240.02 0.52 240.28 5.57 ;
      RECT 239.95 219.01 240.31 219.74 ;
      RECT 240.52 219.01 240.72 219.74 ;
      RECT 240.53 0.3 240.79 5.235 ;
      RECT 241.04 0.52 241.3 7.78 ;
      RECT 241.175 219.01 241.375 219.74 ;
      RECT 241.585 219.01 241.945 219.74 ;
      RECT 241.89 0.52 242.15 4.315 ;
      RECT 242.155 219.01 242.355 219.74 ;
      RECT 242.81 219.01 243.01 219.74 ;
      RECT 243.065 0.52 243.325 2.82 ;
      RECT 243.22 219.01 243.58 219.74 ;
      RECT 243.875 219.01 244.075 219.74 ;
      RECT 244.37 219.01 244.73 219.74 ;
      RECT 245.305 0.18 246.075 0.88 ;
      RECT 245.305 0.18 245.565 12.9 ;
      RECT 245.815 0.18 246.075 12.9 ;
      RECT 244.595 0.52 244.855 2.82 ;
      RECT 244.94 219.01 245.14 219.74 ;
      RECT 246.325 0.155 247.095 0.445 ;
      RECT 246.325 0.155 246.585 13.21 ;
      RECT 246.835 0.155 247.095 13.21 ;
      RECT 245.595 219.01 245.795 219.74 ;
      RECT 246.005 219.01 246.365 219.74 ;
      RECT 246.575 219.01 246.775 219.74 ;
      RECT 247.23 219.01 247.43 219.74 ;
      RECT 247.64 219.01 248 219.74 ;
      RECT 248.295 219.01 248.495 219.74 ;
      RECT 248.79 219.01 249.15 219.74 ;
      RECT 249.03 0.52 249.29 14.115 ;
      RECT 249.36 219.01 249.56 219.74 ;
      RECT 249.54 0.52 249.8 13.45 ;
      RECT 250.015 219.01 250.215 219.74 ;
      RECT 250.56 0.155 251.33 0.445 ;
      RECT 250.56 0.155 250.82 8.665 ;
      RECT 251.07 0.155 251.33 8.665 ;
      RECT 250.05 0.52 250.31 11.315 ;
      RECT 250.425 219.01 250.785 219.74 ;
      RECT 250.995 219.01 251.195 219.74 ;
      RECT 251.58 0.52 251.84 9.955 ;
      RECT 251.65 219.01 251.85 219.74 ;
      RECT 252.06 219.01 252.42 219.74 ;
      RECT 252.715 219.01 252.915 219.74 ;
      RECT 253.21 219.01 253.57 219.74 ;
      RECT 253.62 0.3 253.88 8.7 ;
      RECT 253.78 219.01 253.98 219.74 ;
      RECT 254.435 219.01 254.635 219.74 ;
      RECT 254.13 0.18 254.9 0.88 ;
      RECT 254.845 219.01 255.205 219.74 ;
      RECT 255.415 219.01 255.615 219.74 ;
      RECT 256.07 219.01 256.27 219.74 ;
      RECT 256.325 0.52 256.585 6.28 ;
      RECT 256.48 219.01 256.84 219.74 ;
      RECT 257.135 219.01 257.335 219.74 ;
      RECT 257.7 0.52 257.96 5.57 ;
      RECT 257.63 219.01 257.99 219.74 ;
      RECT 258.2 219.01 258.4 219.74 ;
      RECT 258.21 0.3 258.47 5.235 ;
      RECT 258.72 0.52 258.98 7.78 ;
      RECT 258.855 219.01 259.055 219.74 ;
      RECT 259.265 219.01 259.625 219.74 ;
      RECT 259.835 219.01 260.035 219.74 ;
      RECT 260.66 53.41 260.86 219.74 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 259.24 0 261.17 219.77 ;
      RECT 0 0.52 261.17 219.77 ;
      RECT 258.21 0.3 258.47 219.77 ;
      RECT 256.845 0 257.44 219.77 ;
      RECT 252.1 0 256.065 219.77 ;
      RECT 250.56 0.155 251.33 219.77 ;
      RECT 245.115 0 248.77 219.77 ;
      RECT 243.585 0 244.335 219.77 ;
      RECT 242.41 0 242.805 219.77 ;
      RECT 240.53 0.3 240.79 219.77 ;
      RECT 239.165 0 239.76 219.77 ;
      RECT 234.42 0 238.385 219.77 ;
      RECT 232.88 0.155 233.65 219.77 ;
      RECT 227.435 0 231.09 219.77 ;
      RECT 225.905 0 226.655 219.77 ;
      RECT 224.73 0 225.125 219.77 ;
      RECT 222.85 0.3 223.11 219.77 ;
      RECT 221.485 0 222.08 219.77 ;
      RECT 216.74 0 220.705 219.77 ;
      RECT 215.2 0.155 215.97 219.77 ;
      RECT 209.755 0 213.41 219.77 ;
      RECT 208.225 0 208.975 219.77 ;
      RECT 207.05 0 207.445 219.77 ;
      RECT 205.17 0.3 205.43 219.77 ;
      RECT 203.805 0 204.4 219.77 ;
      RECT 199.06 0 203.025 219.77 ;
      RECT 197.52 0.155 198.29 219.77 ;
      RECT 192.075 0 195.73 219.77 ;
      RECT 190.545 0 191.295 219.77 ;
      RECT 189.37 0 189.765 219.77 ;
      RECT 166.565 0.18 188.59 219.77 ;
      RECT 166.575 0 188.59 219.77 ;
      RECT 161.975 0.3 165.805 219.77 ;
      RECT 158.915 0.18 160.705 219.77 ;
      RECT 153.305 0.3 154.585 219.77 ;
      RECT 150.755 0.3 152.035 219.77 ;
      RECT 149.225 0.3 149.485 219.77 ;
      RECT 146.165 0.3 146.425 219.77 ;
      RECT 144.635 0.3 144.895 219.77 ;
      RECT 136.475 0.3 143.365 219.77 ;
      RECT 126.985 0 134.185 219.77 ;
      RECT 117.805 0.3 124.695 219.77 ;
      RECT 117.815 0 124.695 219.77 ;
      RECT 116.275 0.3 116.535 219.77 ;
      RECT 114.745 0.3 115.005 219.77 ;
      RECT 111.685 0.3 111.945 219.77 ;
      RECT 109.135 0.3 110.415 219.77 ;
      RECT 106.585 0.3 107.865 219.77 ;
      RECT 100.465 0.18 102.255 219.77 ;
      RECT 100.475 0 102.255 219.77 ;
      RECT 95.365 0.3 99.195 219.77 ;
      RECT 72.58 0.18 94.605 219.77 ;
      RECT 71.405 0 71.8 219.77 ;
      RECT 69.875 0 70.625 219.77 ;
      RECT 65.44 0 69.095 219.77 ;
      RECT 62.88 0.155 63.65 219.77 ;
      RECT 58.145 0 62.11 219.77 ;
      RECT 56.77 0 57.365 219.77 ;
      RECT 55.74 0.3 56 219.77 ;
      RECT 53.725 0 54.12 219.77 ;
      RECT 52.195 0 52.945 219.77 ;
      RECT 47.76 0 51.415 219.77 ;
      RECT 45.2 0.155 45.97 219.77 ;
      RECT 40.465 0 44.43 219.77 ;
      RECT 39.09 0 39.685 219.77 ;
      RECT 38.06 0.3 38.32 219.77 ;
      RECT 36.045 0 36.44 219.77 ;
      RECT 34.515 0 35.265 219.77 ;
      RECT 30.08 0 33.735 219.77 ;
      RECT 27.52 0.155 28.29 219.77 ;
      RECT 22.785 0 26.75 219.77 ;
      RECT 21.41 0 22.005 219.77 ;
      RECT 20.38 0.3 20.64 219.77 ;
      RECT 18.365 0 18.76 219.77 ;
      RECT 16.835 0 17.585 219.77 ;
      RECT 12.4 0 16.055 219.77 ;
      RECT 9.84 0.155 10.61 219.77 ;
      RECT 5.105 0 9.07 219.77 ;
      RECT 3.73 0 4.325 219.77 ;
      RECT 2.7 0.3 2.96 219.77 ;
      RECT 0 0 1.93 219.77 ;
      RECT 258.22 0 258.46 219.77 ;
      RECT 240.54 0 240.78 219.77 ;
      RECT 222.86 0 223.1 219.77 ;
      RECT 205.18 0 205.42 219.77 ;
      RECT 161.985 0 165.795 219.77 ;
      RECT 153.315 0 154.575 219.77 ;
      RECT 150.765 0 152.025 219.77 ;
      RECT 149.235 0 149.475 219.77 ;
      RECT 146.175 0 146.415 219.77 ;
      RECT 144.645 0 144.885 219.77 ;
      RECT 136.475 0 143.355 219.77 ;
      RECT 116.285 0 116.525 219.77 ;
      RECT 114.755 0 114.995 219.77 ;
      RECT 111.695 0 111.935 219.77 ;
      RECT 109.145 0 110.405 219.77 ;
      RECT 106.595 0 107.855 219.77 ;
      RECT 95.375 0 99.185 219.77 ;
      RECT 55.75 0 55.99 219.77 ;
      RECT 38.07 0 38.31 219.77 ;
      RECT 20.39 0 20.63 219.77 ;
      RECT 2.71 0 2.95 219.77 ;
      RECT 158.915 0 160.695 219.77 ;
      RECT 72.58 0 94.595 219.77 ;
      RECT 250.57 0 251.32 219.77 ;
      RECT 232.89 0 233.64 219.77 ;
      RECT 215.21 0 215.96 219.77 ;
      RECT 197.53 0 198.28 219.77 ;
      RECT 62.89 0 63.64 219.77 ;
      RECT 45.21 0 45.96 219.77 ;
      RECT 27.53 0 28.28 219.77 ;
      RECT 9.85 0 10.6 219.77 ;
    LAYER Metal3 ;
      RECT 0 0 261.17 219.77 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 170.875 0 188.465 219.77 ;
      RECT 165.725 0 167.545 219.77 ;
      RECT 160.575 0 162.395 219.77 ;
      RECT 255.285 0 261.17 219.77 ;
      RECT 246.445 0 250.345 219.77 ;
      RECT 246.445 47.305 261.17 53.15 ;
      RECT 237.605 0 241.505 219.77 ;
      RECT 228.765 0 232.665 219.77 ;
      RECT 228.765 47.305 241.505 53.15 ;
      RECT 219.925 0 223.825 219.77 ;
      RECT 211.085 0 214.985 219.77 ;
      RECT 211.085 47.305 223.825 53.15 ;
      RECT 202.245 0 206.145 219.77 ;
      RECT 193.405 0 197.305 219.77 ;
      RECT 193.405 47.305 206.145 53.15 ;
      RECT 155.425 0 157.245 219.77 ;
      RECT 150.275 0 152.095 219.77 ;
      RECT 145.125 0 146.945 219.77 ;
      RECT 139.975 0 141.795 219.77 ;
      RECT 134.825 0 136.645 219.77 ;
      RECT 129.675 0 131.495 219.77 ;
      RECT 124.525 0 126.345 219.77 ;
      RECT 119.375 0 121.195 219.77 ;
      RECT 114.225 0 116.045 219.77 ;
      RECT 109.075 0 110.895 219.77 ;
      RECT 103.925 0 105.745 219.77 ;
      RECT 98.775 0 100.595 219.77 ;
      RECT 93.625 0 95.445 219.77 ;
      RECT 72.705 0 90.295 219.77 ;
      RECT 63.865 0 67.765 219.77 ;
      RECT 55.025 0 58.925 219.77 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 219.77 ;
      RECT 37.345 0 41.245 219.77 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 219.77 ;
      RECT 19.665 0 23.565 219.77 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 219.77 ;
      RECT 0 0 5.885 219.77 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_512x8_c2_bm_bist

END LIBRARY
