# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 12:16:39 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_512x16_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_512x16_c2_bm_bist 0 0 ;
  SIZE 236.8 BY 191.34 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 154.57 0 154.83 0.26 ;
    END
  END A_DIN[8]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.97 0 82.23 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.715 0 153.975 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.825 0 83.085 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.73 0 146.99 0.26 ;
    END
  END A_BM[8]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.81 0 90.07 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 148.105 0 148.365 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.435 0 88.695 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 147.24 0 147.5 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.3 0 89.56 0.26 ;
    END
  END A_DOUT[7]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 224.11 0 226.92 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.87 0 215.68 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 201.63 0 204.44 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.39 0 193.2 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.15 0 181.96 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.91 0 170.72 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.67 0 159.48 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.43 0 148.24 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.02 0 137.83 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.72 0 127.53 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.27 0 112.08 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 98.97 0 101.78 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 191.34 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 0 232.54 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 0 221.3 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 0 210.06 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 0 198.82 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 0 187.58 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 0 176.34 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 0 165.1 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 0 153.86 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.87 0 132.68 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.57 0 122.38 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.42 0 117.23 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 104.12 0 106.93 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 38.825 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 45.465 232.54 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 45.465 221.3 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 45.465 210.06 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 45.465 198.82 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 45.465 187.58 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 45.465 176.34 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 45.465 165.1 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 45.465 153.86 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 45.465 85.75 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 45.465 74.51 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 45.465 63.27 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 45.465 52.03 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 45.465 40.79 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 45.465 29.55 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 45.465 18.31 191.34 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 45.465 7.07 191.34 ;
    END
  END VDDARRAY!
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 165.81 0 166.07 0.26 ;
    END
  END A_DIN[9]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.73 0 70.99 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 164.955 0 165.215 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 71.585 0 71.845 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.97 0 158.23 0.26 ;
    END
  END A_BM[9]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.57 0 78.83 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 159.345 0 159.605 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.195 0 77.455 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.48 0 158.74 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.06 0 78.32 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 177.05 0 177.31 0.26 ;
    END
  END A_DIN[10]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 59.49 0 59.75 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.195 0 176.455 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.345 0 60.605 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 169.21 0 169.47 0.26 ;
    END
  END A_BM[10]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.33 0 67.59 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 170.585 0 170.845 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 65.955 0 66.215 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 169.72 0 169.98 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.82 0 67.08 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.29 0 188.55 0.26 ;
    END
  END A_DIN[11]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 48.25 0 48.51 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 187.435 0 187.695 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 49.105 0 49.365 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 180.45 0 180.71 0.26 ;
    END
  END A_BM[11]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.09 0 56.35 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.825 0 182.085 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.715 0 54.975 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 180.96 0 181.22 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.58 0 55.84 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 199.53 0 199.79 0.26 ;
    END
  END A_DIN[12]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.01 0 37.27 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 198.675 0 198.935 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.865 0 38.125 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 191.69 0 191.95 0.26 ;
    END
  END A_BM[12]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.85 0 45.11 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.065 0 193.325 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 43.475 0 43.735 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.2 0 192.46 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.34 0 44.6 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 210.77 0 211.03 0.26 ;
    END
  END A_DIN[13]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 25.77 0 26.03 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 209.915 0 210.175 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 26.625 0 26.885 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.93 0 203.19 0.26 ;
    END
  END A_BM[13]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.61 0 33.87 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.305 0 204.565 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.235 0 32.495 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.44 0 203.7 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.1 0 33.36 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 222.01 0 222.27 0.26 ;
    END
  END A_DIN[14]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.53 0 14.79 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221.155 0 221.415 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.385 0 15.645 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.17 0 214.43 0.26 ;
    END
  END A_BM[14]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.37 0 22.63 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.545 0 215.805 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.995 0 21.255 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.68 0 214.94 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 21.86 0 22.12 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 233.25 0 233.51 0.26 ;
    END
  END A_DIN[15]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.29 0 3.55 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.395 0 232.655 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.145 0 4.405 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 225.41 0 225.67 0.26 ;
    END
  END A_BM[15]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.13 0 11.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.785 0 227.045 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.755 0 10.015 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 225.92 0 226.18 0.26 ;
    END
  END A_DOUT[15]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.62 0 10.88 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 45.223301 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.6 0 114.86 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.184466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.19 0 119.45 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 39.656958 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.09 0 114.35 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.618123 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 118.68 0 118.94 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.25 0 122.51 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.76 0 123.02 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.23 0 121.49 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.74 0 122 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.63754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.8 0 125.06 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.317152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.29 0 124.55 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 70.245955 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.78 0 124.04 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 68.925566 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.27 0 123.53 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 55.436893 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.36 0 102.62 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 54.065721 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.87 0 103.13 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 62.724919 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.38 0 103.64 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.404531 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.89 0 104.15 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.740105 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 132.45 0 132.71 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.204381 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 132.96 0 133.22 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.56 0 112.82 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.796863 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.13 0 116.39 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.62 0 115.88 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.07 0 113.33 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 18.532819 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.49 0 134.75 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 114.62575 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 16.0875 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.213636 LAYER Metal2 ;
      ANTENNAMAXAREACAR 17.397871 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.11 0 115.37 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.03 0 111.29 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.66 0 117.92 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.15 0 117.41 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.54 0 111.8 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 236.8 191.34 ;
    LAYER Metal2 ;
      RECT 0.105 45.465 0.305 191.315 ;
      RECT 1.1 190.585 1.3 191.315 ;
      RECT 3.29 0.52 3.55 5.16 ;
      RECT 2.77 4.9 3.55 5.16 ;
      RECT 2.77 4.9 3.03 6.64 ;
      RECT 1.92 190.585 2.12 191.315 ;
      RECT 2.415 190.585 2.615 191.315 ;
      RECT 2.915 190.585 3.115 191.315 ;
      RECT 3.415 190.585 3.615 191.315 ;
      RECT 3.91 190.585 4.11 191.315 ;
      RECT 4.655 0.17 5.425 0.94 ;
      RECT 4.655 0.17 4.915 12.9 ;
      RECT 5.165 0.17 5.425 12.9 ;
      RECT 4.145 0.52 4.405 5.815 ;
      RECT 4.73 190.585 4.93 191.315 ;
      RECT 5.675 0.17 6.445 0.43 ;
      RECT 5.675 0.17 5.935 11.5 ;
      RECT 6.185 0.17 6.445 11.5 ;
      RECT 5.225 190.585 5.425 191.315 ;
      RECT 5.725 190.585 5.925 191.315 ;
      RECT 6.225 190.585 6.425 191.315 ;
      RECT 7.715 0.17 8.485 0.43 ;
      RECT 7.715 0.17 7.975 10.48 ;
      RECT 8.225 0.17 8.485 10.99 ;
      RECT 6.72 190.585 6.92 191.315 ;
      RECT 7.54 190.585 7.74 191.315 ;
      RECT 8.735 0.17 9.505 0.94 ;
      RECT 8.735 0.17 8.995 8.7 ;
      RECT 9.245 0.17 9.505 12.9 ;
      RECT 8.035 190.585 8.235 191.315 ;
      RECT 8.535 190.585 8.735 191.315 ;
      RECT 9.035 190.585 9.235 191.315 ;
      RECT 9.53 190.585 9.73 191.315 ;
      RECT 9.755 0.52 10.015 2.485 ;
      RECT 10.35 190.585 10.55 191.315 ;
      RECT 10.62 0.52 10.88 14.11 ;
      RECT 10.845 190.585 11.045 191.315 ;
      RECT 11.13 0.52 11.39 2.335 ;
      RECT 11.345 190.585 11.545 191.315 ;
      RECT 11.845 190.585 12.045 191.315 ;
      RECT 12.34 190.585 12.54 191.315 ;
      RECT 14.53 0.52 14.79 5.16 ;
      RECT 14.01 4.9 14.79 5.16 ;
      RECT 14.01 4.9 14.27 6.64 ;
      RECT 13.16 190.585 13.36 191.315 ;
      RECT 13.655 190.585 13.855 191.315 ;
      RECT 14.155 190.585 14.355 191.315 ;
      RECT 14.655 190.585 14.855 191.315 ;
      RECT 15.15 190.585 15.35 191.315 ;
      RECT 15.895 0.17 16.665 0.94 ;
      RECT 15.895 0.17 16.155 12.9 ;
      RECT 16.405 0.17 16.665 12.9 ;
      RECT 15.385 0.52 15.645 5.815 ;
      RECT 15.97 190.585 16.17 191.315 ;
      RECT 16.915 0.17 17.685 0.43 ;
      RECT 16.915 0.17 17.175 11.5 ;
      RECT 17.425 0.17 17.685 11.5 ;
      RECT 16.465 190.585 16.665 191.315 ;
      RECT 16.965 190.585 17.165 191.315 ;
      RECT 17.465 190.585 17.665 191.315 ;
      RECT 18.955 0.17 19.725 0.43 ;
      RECT 18.955 0.17 19.215 10.48 ;
      RECT 19.465 0.17 19.725 10.99 ;
      RECT 17.96 190.585 18.16 191.315 ;
      RECT 18.78 190.585 18.98 191.315 ;
      RECT 19.975 0.17 20.745 0.94 ;
      RECT 19.975 0.17 20.235 8.7 ;
      RECT 20.485 0.17 20.745 12.9 ;
      RECT 19.275 190.585 19.475 191.315 ;
      RECT 19.775 190.585 19.975 191.315 ;
      RECT 20.275 190.585 20.475 191.315 ;
      RECT 20.77 190.585 20.97 191.315 ;
      RECT 20.995 0.52 21.255 2.485 ;
      RECT 21.59 190.585 21.79 191.315 ;
      RECT 21.86 0.52 22.12 14.11 ;
      RECT 22.085 190.585 22.285 191.315 ;
      RECT 22.37 0.52 22.63 2.335 ;
      RECT 22.585 190.585 22.785 191.315 ;
      RECT 23.085 190.585 23.285 191.315 ;
      RECT 23.58 190.585 23.78 191.315 ;
      RECT 25.77 0.52 26.03 5.16 ;
      RECT 25.25 4.9 26.03 5.16 ;
      RECT 25.25 4.9 25.51 6.64 ;
      RECT 24.4 190.585 24.6 191.315 ;
      RECT 24.895 190.585 25.095 191.315 ;
      RECT 25.395 190.585 25.595 191.315 ;
      RECT 25.895 190.585 26.095 191.315 ;
      RECT 26.39 190.585 26.59 191.315 ;
      RECT 27.135 0.17 27.905 0.94 ;
      RECT 27.135 0.17 27.395 12.9 ;
      RECT 27.645 0.17 27.905 12.9 ;
      RECT 26.625 0.52 26.885 5.815 ;
      RECT 27.21 190.585 27.41 191.315 ;
      RECT 28.155 0.17 28.925 0.43 ;
      RECT 28.155 0.17 28.415 11.5 ;
      RECT 28.665 0.17 28.925 11.5 ;
      RECT 27.705 190.585 27.905 191.315 ;
      RECT 28.205 190.585 28.405 191.315 ;
      RECT 28.705 190.585 28.905 191.315 ;
      RECT 30.195 0.17 30.965 0.43 ;
      RECT 30.195 0.17 30.455 10.48 ;
      RECT 30.705 0.17 30.965 10.99 ;
      RECT 29.2 190.585 29.4 191.315 ;
      RECT 30.02 190.585 30.22 191.315 ;
      RECT 31.215 0.17 31.985 0.94 ;
      RECT 31.215 0.17 31.475 8.7 ;
      RECT 31.725 0.17 31.985 12.9 ;
      RECT 30.515 190.585 30.715 191.315 ;
      RECT 31.015 190.585 31.215 191.315 ;
      RECT 31.515 190.585 31.715 191.315 ;
      RECT 32.01 190.585 32.21 191.315 ;
      RECT 32.235 0.52 32.495 2.485 ;
      RECT 32.83 190.585 33.03 191.315 ;
      RECT 33.1 0.52 33.36 14.11 ;
      RECT 33.325 190.585 33.525 191.315 ;
      RECT 33.61 0.52 33.87 2.335 ;
      RECT 33.825 190.585 34.025 191.315 ;
      RECT 34.325 190.585 34.525 191.315 ;
      RECT 34.82 190.585 35.02 191.315 ;
      RECT 37.01 0.52 37.27 5.16 ;
      RECT 36.49 4.9 37.27 5.16 ;
      RECT 36.49 4.9 36.75 6.64 ;
      RECT 35.64 190.585 35.84 191.315 ;
      RECT 36.135 190.585 36.335 191.315 ;
      RECT 36.635 190.585 36.835 191.315 ;
      RECT 37.135 190.585 37.335 191.315 ;
      RECT 37.63 190.585 37.83 191.315 ;
      RECT 38.375 0.17 39.145 0.94 ;
      RECT 38.375 0.17 38.635 12.9 ;
      RECT 38.885 0.17 39.145 12.9 ;
      RECT 37.865 0.52 38.125 5.815 ;
      RECT 38.45 190.585 38.65 191.315 ;
      RECT 39.395 0.17 40.165 0.43 ;
      RECT 39.395 0.17 39.655 11.5 ;
      RECT 39.905 0.17 40.165 11.5 ;
      RECT 38.945 190.585 39.145 191.315 ;
      RECT 39.445 190.585 39.645 191.315 ;
      RECT 39.945 190.585 40.145 191.315 ;
      RECT 41.435 0.17 42.205 0.43 ;
      RECT 41.435 0.17 41.695 10.48 ;
      RECT 41.945 0.17 42.205 10.99 ;
      RECT 40.44 190.585 40.64 191.315 ;
      RECT 41.26 190.585 41.46 191.315 ;
      RECT 42.455 0.17 43.225 0.94 ;
      RECT 42.455 0.17 42.715 8.7 ;
      RECT 42.965 0.17 43.225 12.9 ;
      RECT 41.755 190.585 41.955 191.315 ;
      RECT 42.255 190.585 42.455 191.315 ;
      RECT 42.755 190.585 42.955 191.315 ;
      RECT 43.25 190.585 43.45 191.315 ;
      RECT 43.475 0.52 43.735 2.485 ;
      RECT 44.07 190.585 44.27 191.315 ;
      RECT 44.34 0.52 44.6 14.11 ;
      RECT 44.565 190.585 44.765 191.315 ;
      RECT 44.85 0.52 45.11 2.335 ;
      RECT 45.065 190.585 45.265 191.315 ;
      RECT 45.565 190.585 45.765 191.315 ;
      RECT 46.06 190.585 46.26 191.315 ;
      RECT 48.25 0.52 48.51 5.16 ;
      RECT 47.73 4.9 48.51 5.16 ;
      RECT 47.73 4.9 47.99 6.64 ;
      RECT 46.88 190.585 47.08 191.315 ;
      RECT 47.375 190.585 47.575 191.315 ;
      RECT 47.875 190.585 48.075 191.315 ;
      RECT 48.375 190.585 48.575 191.315 ;
      RECT 48.87 190.585 49.07 191.315 ;
      RECT 49.615 0.17 50.385 0.94 ;
      RECT 49.615 0.17 49.875 12.9 ;
      RECT 50.125 0.17 50.385 12.9 ;
      RECT 49.105 0.52 49.365 5.815 ;
      RECT 49.69 190.585 49.89 191.315 ;
      RECT 50.635 0.17 51.405 0.43 ;
      RECT 50.635 0.17 50.895 11.5 ;
      RECT 51.145 0.17 51.405 11.5 ;
      RECT 50.185 190.585 50.385 191.315 ;
      RECT 50.685 190.585 50.885 191.315 ;
      RECT 51.185 190.585 51.385 191.315 ;
      RECT 52.675 0.17 53.445 0.43 ;
      RECT 52.675 0.17 52.935 10.48 ;
      RECT 53.185 0.17 53.445 10.99 ;
      RECT 51.68 190.585 51.88 191.315 ;
      RECT 52.5 190.585 52.7 191.315 ;
      RECT 53.695 0.17 54.465 0.94 ;
      RECT 53.695 0.17 53.955 8.7 ;
      RECT 54.205 0.17 54.465 12.9 ;
      RECT 52.995 190.585 53.195 191.315 ;
      RECT 53.495 190.585 53.695 191.315 ;
      RECT 53.995 190.585 54.195 191.315 ;
      RECT 54.49 190.585 54.69 191.315 ;
      RECT 54.715 0.52 54.975 2.485 ;
      RECT 55.31 190.585 55.51 191.315 ;
      RECT 55.58 0.52 55.84 14.11 ;
      RECT 55.805 190.585 56.005 191.315 ;
      RECT 56.09 0.52 56.35 2.335 ;
      RECT 56.305 190.585 56.505 191.315 ;
      RECT 56.805 190.585 57.005 191.315 ;
      RECT 57.3 190.585 57.5 191.315 ;
      RECT 59.49 0.52 59.75 5.16 ;
      RECT 58.97 4.9 59.75 5.16 ;
      RECT 58.97 4.9 59.23 6.64 ;
      RECT 58.12 190.585 58.32 191.315 ;
      RECT 58.615 190.585 58.815 191.315 ;
      RECT 59.115 190.585 59.315 191.315 ;
      RECT 59.615 190.585 59.815 191.315 ;
      RECT 60.11 190.585 60.31 191.315 ;
      RECT 60.855 0.17 61.625 0.94 ;
      RECT 60.855 0.17 61.115 12.9 ;
      RECT 61.365 0.17 61.625 12.9 ;
      RECT 60.345 0.52 60.605 5.815 ;
      RECT 60.93 190.585 61.13 191.315 ;
      RECT 61.875 0.17 62.645 0.43 ;
      RECT 61.875 0.17 62.135 11.5 ;
      RECT 62.385 0.17 62.645 11.5 ;
      RECT 61.425 190.585 61.625 191.315 ;
      RECT 61.925 190.585 62.125 191.315 ;
      RECT 62.425 190.585 62.625 191.315 ;
      RECT 63.915 0.17 64.685 0.43 ;
      RECT 63.915 0.17 64.175 10.48 ;
      RECT 64.425 0.17 64.685 10.99 ;
      RECT 62.92 190.585 63.12 191.315 ;
      RECT 63.74 190.585 63.94 191.315 ;
      RECT 64.935 0.17 65.705 0.94 ;
      RECT 64.935 0.17 65.195 8.7 ;
      RECT 65.445 0.17 65.705 12.9 ;
      RECT 64.235 190.585 64.435 191.315 ;
      RECT 64.735 190.585 64.935 191.315 ;
      RECT 65.235 190.585 65.435 191.315 ;
      RECT 65.73 190.585 65.93 191.315 ;
      RECT 65.955 0.52 66.215 2.485 ;
      RECT 66.55 190.585 66.75 191.315 ;
      RECT 66.82 0.52 67.08 14.11 ;
      RECT 67.045 190.585 67.245 191.315 ;
      RECT 67.33 0.52 67.59 2.335 ;
      RECT 67.545 190.585 67.745 191.315 ;
      RECT 68.045 190.585 68.245 191.315 ;
      RECT 68.54 190.585 68.74 191.315 ;
      RECT 70.73 0.52 70.99 5.16 ;
      RECT 70.21 4.9 70.99 5.16 ;
      RECT 70.21 4.9 70.47 6.64 ;
      RECT 69.36 190.585 69.56 191.315 ;
      RECT 69.855 190.585 70.055 191.315 ;
      RECT 70.355 190.585 70.555 191.315 ;
      RECT 70.855 190.585 71.055 191.315 ;
      RECT 71.35 190.585 71.55 191.315 ;
      RECT 72.095 0.17 72.865 0.94 ;
      RECT 72.095 0.17 72.355 12.9 ;
      RECT 72.605 0.17 72.865 12.9 ;
      RECT 71.585 0.52 71.845 5.815 ;
      RECT 72.17 190.585 72.37 191.315 ;
      RECT 73.115 0.17 73.885 0.43 ;
      RECT 73.115 0.17 73.375 11.5 ;
      RECT 73.625 0.17 73.885 11.5 ;
      RECT 72.665 190.585 72.865 191.315 ;
      RECT 73.165 190.585 73.365 191.315 ;
      RECT 73.665 190.585 73.865 191.315 ;
      RECT 75.155 0.17 75.925 0.43 ;
      RECT 75.155 0.17 75.415 10.48 ;
      RECT 75.665 0.17 75.925 10.99 ;
      RECT 74.16 190.585 74.36 191.315 ;
      RECT 74.98 190.585 75.18 191.315 ;
      RECT 76.175 0.17 76.945 0.94 ;
      RECT 76.175 0.17 76.435 8.7 ;
      RECT 76.685 0.17 76.945 12.9 ;
      RECT 75.475 190.585 75.675 191.315 ;
      RECT 75.975 190.585 76.175 191.315 ;
      RECT 76.475 190.585 76.675 191.315 ;
      RECT 76.97 190.585 77.17 191.315 ;
      RECT 77.195 0.52 77.455 2.485 ;
      RECT 77.79 190.585 77.99 191.315 ;
      RECT 78.06 0.52 78.32 14.11 ;
      RECT 78.285 190.585 78.485 191.315 ;
      RECT 78.57 0.52 78.83 2.335 ;
      RECT 78.785 190.585 78.985 191.315 ;
      RECT 79.285 190.585 79.485 191.315 ;
      RECT 79.78 190.585 79.98 191.315 ;
      RECT 81.97 0.52 82.23 5.16 ;
      RECT 81.45 4.9 82.23 5.16 ;
      RECT 81.45 4.9 81.71 6.64 ;
      RECT 80.6 190.585 80.8 191.315 ;
      RECT 81.095 190.585 81.295 191.315 ;
      RECT 81.595 190.585 81.795 191.315 ;
      RECT 82.095 190.585 82.295 191.315 ;
      RECT 82.59 190.585 82.79 191.315 ;
      RECT 83.335 0.17 84.105 0.94 ;
      RECT 83.335 0.17 83.595 12.9 ;
      RECT 83.845 0.17 84.105 12.9 ;
      RECT 82.825 0.52 83.085 5.815 ;
      RECT 83.41 190.585 83.61 191.315 ;
      RECT 84.355 0.17 85.125 0.43 ;
      RECT 84.355 0.17 84.615 11.5 ;
      RECT 84.865 0.17 85.125 11.5 ;
      RECT 83.905 190.585 84.105 191.315 ;
      RECT 84.405 190.585 84.605 191.315 ;
      RECT 84.905 190.585 85.105 191.315 ;
      RECT 86.395 0.17 87.165 0.43 ;
      RECT 86.395 0.17 86.655 10.48 ;
      RECT 86.905 0.17 87.165 10.99 ;
      RECT 85.4 190.585 85.6 191.315 ;
      RECT 86.22 190.585 86.42 191.315 ;
      RECT 87.415 0.17 88.185 0.94 ;
      RECT 87.415 0.17 87.675 8.7 ;
      RECT 87.925 0.17 88.185 12.9 ;
      RECT 86.715 190.585 86.915 191.315 ;
      RECT 87.215 190.585 87.415 191.315 ;
      RECT 87.715 190.585 87.915 191.315 ;
      RECT 88.21 190.585 88.41 191.315 ;
      RECT 88.435 0.52 88.695 2.485 ;
      RECT 89.03 190.585 89.23 191.315 ;
      RECT 89.3 0.52 89.56 14.11 ;
      RECT 89.525 190.585 89.725 191.315 ;
      RECT 89.81 0.52 90.07 2.335 ;
      RECT 90.025 190.585 90.225 191.315 ;
      RECT 90.525 190.585 90.725 191.315 ;
      RECT 92.515 0.17 93.285 0.43 ;
      RECT 92.515 0.17 92.775 8.7 ;
      RECT 93.025 0.17 93.285 8.7 ;
      RECT 93.535 0.17 94.305 0.94 ;
      RECT 93.535 0.17 93.795 8.7 ;
      RECT 94.045 0.17 94.305 8.7 ;
      RECT 94.555 0.17 95.325 0.43 ;
      RECT 94.555 0.17 94.815 8.7 ;
      RECT 95.065 0.17 95.325 8.7 ;
      RECT 95.575 0.17 96.345 0.94 ;
      RECT 95.575 0.17 95.835 8.7 ;
      RECT 96.085 0.17 96.345 8.7 ;
      RECT 96.595 0.17 97.365 0.43 ;
      RECT 96.595 0.17 96.855 8.7 ;
      RECT 97.105 0.17 97.365 8.7 ;
      RECT 97.615 0.17 98.385 0.94 ;
      RECT 97.615 0.17 97.875 8.7 ;
      RECT 98.125 0.17 98.385 8.7 ;
      RECT 91.02 190.585 91.22 191.315 ;
      RECT 91.84 190.585 92.04 191.315 ;
      RECT 92.835 190.585 93.035 191.315 ;
      RECT 100.32 0.17 101.09 0.94 ;
      RECT 100.32 0.17 100.58 8.7 ;
      RECT 100.83 0.17 101.09 8.7 ;
      RECT 98.79 0.3 99.05 8.7 ;
      RECT 99.3 0 99.56 8.7 ;
      RECT 99.81 0 100.07 8.7 ;
      RECT 101.34 0 101.6 8.7 ;
      RECT 101.85 0 102.11 8.7 ;
      RECT 102.36 0.52 102.62 8.7 ;
      RECT 102.87 0.52 103.13 8.7 ;
      RECT 103.38 0.52 103.64 8.7 ;
      RECT 105.42 0.17 106.19 0.94 ;
      RECT 105.42 0.17 105.68 8.7 ;
      RECT 105.93 0.17 106.19 8.7 ;
      RECT 106.44 0.17 107.21 0.43 ;
      RECT 106.44 0.17 106.7 8.7 ;
      RECT 106.95 0.17 107.21 8.7 ;
      RECT 103.89 0.52 104.15 8.7 ;
      RECT 104.4 0 104.66 8.7 ;
      RECT 104.91 0 105.17 8.7 ;
      RECT 107.46 0.3 107.72 8.7 ;
      RECT 107.97 0.3 108.23 8.7 ;
      RECT 110.01 0.17 110.78 0.94 ;
      RECT 110.01 0.17 110.27 8.7 ;
      RECT 110.52 0.17 110.78 8.7 ;
      RECT 108.48 0.3 108.74 8.7 ;
      RECT 108.99 0.3 109.25 8.7 ;
      RECT 109.5 0.3 109.76 8.7 ;
      RECT 111.03 0.52 111.29 8.7 ;
      RECT 111.54 0.52 111.8 8.7 ;
      RECT 112.05 0.3 112.31 8.7 ;
      RECT 112.56 0.52 112.82 8.7 ;
      RECT 113.07 0.52 113.33 8.7 ;
      RECT 113.58 0.3 113.84 8.7 ;
      RECT 114.09 0.52 114.35 8.7 ;
      RECT 114.6 0.52 114.86 8.7 ;
      RECT 115.11 0.52 115.37 8.7 ;
      RECT 115.62 0.52 115.88 8.7 ;
      RECT 116.13 0.52 116.39 8.7 ;
      RECT 116.64 0.3 116.9 8.7 ;
      RECT 117.15 0.52 117.41 8.7 ;
      RECT 117.66 0.52 117.92 8.7 ;
      RECT 118.17 0.3 118.43 8.7 ;
      RECT 120.21 0.17 120.98 0.94 ;
      RECT 120.21 0.17 120.47 8.7 ;
      RECT 120.72 0.17 120.98 8.7 ;
      RECT 118.68 0.52 118.94 8.7 ;
      RECT 119.19 0.52 119.45 8.7 ;
      RECT 119.7 0.3 119.96 8.7 ;
      RECT 121.23 0.52 121.49 8.7 ;
      RECT 121.74 0.52 122 8.7 ;
      RECT 122.25 0.52 122.51 8.7 ;
      RECT 122.76 0.52 123.02 8.7 ;
      RECT 123.27 0.52 123.53 8.7 ;
      RECT 123.78 0.52 124.04 8.7 ;
      RECT 124.29 0.52 124.55 8.7 ;
      RECT 126.33 0.17 127.1 0.94 ;
      RECT 126.33 0.17 126.59 8.7 ;
      RECT 126.84 0.17 127.1 8.7 ;
      RECT 124.8 0.52 125.06 8.7 ;
      RECT 125.31 0 125.57 8.7 ;
      RECT 125.82 0 126.08 8.7 ;
      RECT 127.35 0 127.61 8.7 ;
      RECT 129.39 0.17 130.16 0.43 ;
      RECT 129.39 0.17 129.65 8.7 ;
      RECT 129.9 0.17 130.16 8.7 ;
      RECT 127.86 0 128.12 8.7 ;
      RECT 128.37 0.3 128.63 8.7 ;
      RECT 128.88 0.3 129.14 8.7 ;
      RECT 130.41 0.3 130.67 8.7 ;
      RECT 130.92 0.3 131.18 8.7 ;
      RECT 131.43 0.3 131.69 8.7 ;
      RECT 131.94 0.3 132.2 8.7 ;
      RECT 132.45 0.52 132.71 8.7 ;
      RECT 132.96 0.52 133.22 8.7 ;
      RECT 135 0.17 135.77 0.43 ;
      RECT 135 0.17 135.26 8.7 ;
      RECT 135.51 0.17 135.77 8.7 ;
      RECT 136.02 0.17 136.79 0.94 ;
      RECT 136.02 0.17 136.28 25.5 ;
      RECT 136.53 0.17 136.79 33.9 ;
      RECT 137.04 0.17 137.81 0.43 ;
      RECT 137.04 0.17 137.3 8.7 ;
      RECT 137.55 0.17 137.81 8.7 ;
      RECT 138.415 0.17 139.185 0.94 ;
      RECT 138.415 0.17 138.675 8.7 ;
      RECT 138.925 0.17 139.185 8.7 ;
      RECT 139.435 0.17 140.205 0.43 ;
      RECT 139.435 0.17 139.695 8.7 ;
      RECT 139.945 0.17 140.205 8.7 ;
      RECT 140.455 0.17 141.225 0.94 ;
      RECT 140.455 0.17 140.715 8.7 ;
      RECT 140.965 0.17 141.225 8.7 ;
      RECT 141.475 0.17 142.245 0.43 ;
      RECT 141.475 0.17 141.735 8.7 ;
      RECT 141.985 0.17 142.245 8.7 ;
      RECT 142.495 0.17 143.265 0.94 ;
      RECT 142.495 0.17 142.755 8.7 ;
      RECT 143.005 0.17 143.265 8.7 ;
      RECT 133.47 0.3 133.73 8.7 ;
      RECT 143.515 0.17 144.285 0.43 ;
      RECT 143.515 0.17 143.775 8.7 ;
      RECT 144.025 0.17 144.285 8.7 ;
      RECT 133.98 0.3 134.24 8.7 ;
      RECT 134.49 0.52 134.75 8.7 ;
      RECT 143.765 190.585 143.965 191.315 ;
      RECT 144.76 190.585 144.96 191.315 ;
      RECT 145.58 190.585 145.78 191.315 ;
      RECT 146.075 190.585 146.275 191.315 ;
      RECT 146.575 190.585 146.775 191.315 ;
      RECT 146.73 0.52 146.99 2.335 ;
      RECT 147.075 190.585 147.275 191.315 ;
      RECT 147.24 0.52 147.5 14.11 ;
      RECT 147.57 190.585 147.77 191.315 ;
      RECT 148.615 0.17 149.385 0.94 ;
      RECT 149.125 0.17 149.385 8.7 ;
      RECT 148.615 0.17 148.875 12.9 ;
      RECT 148.105 0.52 148.365 2.485 ;
      RECT 148.39 190.585 148.59 191.315 ;
      RECT 149.635 0.17 150.405 0.43 ;
      RECT 150.145 0.17 150.405 10.48 ;
      RECT 149.635 0.17 149.895 10.99 ;
      RECT 148.885 190.585 149.085 191.315 ;
      RECT 149.385 190.585 149.585 191.315 ;
      RECT 149.885 190.585 150.085 191.315 ;
      RECT 150.38 190.585 150.58 191.315 ;
      RECT 151.675 0.17 152.445 0.43 ;
      RECT 151.675 0.17 151.935 11.5 ;
      RECT 152.185 0.17 152.445 11.5 ;
      RECT 151.2 190.585 151.4 191.315 ;
      RECT 151.695 190.585 151.895 191.315 ;
      RECT 152.695 0.17 153.465 0.94 ;
      RECT 152.695 0.17 152.955 12.9 ;
      RECT 153.205 0.17 153.465 12.9 ;
      RECT 152.195 190.585 152.395 191.315 ;
      RECT 152.695 190.585 152.895 191.315 ;
      RECT 153.19 190.585 153.39 191.315 ;
      RECT 153.715 0.52 153.975 5.815 ;
      RECT 154.57 0.52 154.83 5.16 ;
      RECT 154.57 4.9 155.35 5.16 ;
      RECT 155.09 4.9 155.35 6.64 ;
      RECT 154.01 190.585 154.21 191.315 ;
      RECT 154.505 190.585 154.705 191.315 ;
      RECT 155.005 190.585 155.205 191.315 ;
      RECT 155.505 190.585 155.705 191.315 ;
      RECT 156 190.585 156.2 191.315 ;
      RECT 156.82 190.585 157.02 191.315 ;
      RECT 157.315 190.585 157.515 191.315 ;
      RECT 157.815 190.585 158.015 191.315 ;
      RECT 157.97 0.52 158.23 2.335 ;
      RECT 158.315 190.585 158.515 191.315 ;
      RECT 158.48 0.52 158.74 14.11 ;
      RECT 158.81 190.585 159.01 191.315 ;
      RECT 159.855 0.17 160.625 0.94 ;
      RECT 160.365 0.17 160.625 8.7 ;
      RECT 159.855 0.17 160.115 12.9 ;
      RECT 159.345 0.52 159.605 2.485 ;
      RECT 159.63 190.585 159.83 191.315 ;
      RECT 160.875 0.17 161.645 0.43 ;
      RECT 161.385 0.17 161.645 10.48 ;
      RECT 160.875 0.17 161.135 10.99 ;
      RECT 160.125 190.585 160.325 191.315 ;
      RECT 160.625 190.585 160.825 191.315 ;
      RECT 161.125 190.585 161.325 191.315 ;
      RECT 161.62 190.585 161.82 191.315 ;
      RECT 162.915 0.17 163.685 0.43 ;
      RECT 162.915 0.17 163.175 11.5 ;
      RECT 163.425 0.17 163.685 11.5 ;
      RECT 162.44 190.585 162.64 191.315 ;
      RECT 162.935 190.585 163.135 191.315 ;
      RECT 163.935 0.17 164.705 0.94 ;
      RECT 163.935 0.17 164.195 12.9 ;
      RECT 164.445 0.17 164.705 12.9 ;
      RECT 163.435 190.585 163.635 191.315 ;
      RECT 163.935 190.585 164.135 191.315 ;
      RECT 164.43 190.585 164.63 191.315 ;
      RECT 164.955 0.52 165.215 5.815 ;
      RECT 165.81 0.52 166.07 5.16 ;
      RECT 165.81 4.9 166.59 5.16 ;
      RECT 166.33 4.9 166.59 6.64 ;
      RECT 165.25 190.585 165.45 191.315 ;
      RECT 165.745 190.585 165.945 191.315 ;
      RECT 166.245 190.585 166.445 191.315 ;
      RECT 166.745 190.585 166.945 191.315 ;
      RECT 167.24 190.585 167.44 191.315 ;
      RECT 168.06 190.585 168.26 191.315 ;
      RECT 168.555 190.585 168.755 191.315 ;
      RECT 169.055 190.585 169.255 191.315 ;
      RECT 169.21 0.52 169.47 2.335 ;
      RECT 169.555 190.585 169.755 191.315 ;
      RECT 169.72 0.52 169.98 14.11 ;
      RECT 170.05 190.585 170.25 191.315 ;
      RECT 171.095 0.17 171.865 0.94 ;
      RECT 171.605 0.17 171.865 8.7 ;
      RECT 171.095 0.17 171.355 12.9 ;
      RECT 170.585 0.52 170.845 2.485 ;
      RECT 170.87 190.585 171.07 191.315 ;
      RECT 172.115 0.17 172.885 0.43 ;
      RECT 172.625 0.17 172.885 10.48 ;
      RECT 172.115 0.17 172.375 10.99 ;
      RECT 171.365 190.585 171.565 191.315 ;
      RECT 171.865 190.585 172.065 191.315 ;
      RECT 172.365 190.585 172.565 191.315 ;
      RECT 172.86 190.585 173.06 191.315 ;
      RECT 174.155 0.17 174.925 0.43 ;
      RECT 174.155 0.17 174.415 11.5 ;
      RECT 174.665 0.17 174.925 11.5 ;
      RECT 173.68 190.585 173.88 191.315 ;
      RECT 174.175 190.585 174.375 191.315 ;
      RECT 175.175 0.17 175.945 0.94 ;
      RECT 175.175 0.17 175.435 12.9 ;
      RECT 175.685 0.17 175.945 12.9 ;
      RECT 174.675 190.585 174.875 191.315 ;
      RECT 175.175 190.585 175.375 191.315 ;
      RECT 175.67 190.585 175.87 191.315 ;
      RECT 176.195 0.52 176.455 5.815 ;
      RECT 177.05 0.52 177.31 5.16 ;
      RECT 177.05 4.9 177.83 5.16 ;
      RECT 177.57 4.9 177.83 6.64 ;
      RECT 176.49 190.585 176.69 191.315 ;
      RECT 176.985 190.585 177.185 191.315 ;
      RECT 177.485 190.585 177.685 191.315 ;
      RECT 177.985 190.585 178.185 191.315 ;
      RECT 178.48 190.585 178.68 191.315 ;
      RECT 179.3 190.585 179.5 191.315 ;
      RECT 179.795 190.585 179.995 191.315 ;
      RECT 180.295 190.585 180.495 191.315 ;
      RECT 180.45 0.52 180.71 2.335 ;
      RECT 180.795 190.585 180.995 191.315 ;
      RECT 180.96 0.52 181.22 14.11 ;
      RECT 181.29 190.585 181.49 191.315 ;
      RECT 182.335 0.17 183.105 0.94 ;
      RECT 182.845 0.17 183.105 8.7 ;
      RECT 182.335 0.17 182.595 12.9 ;
      RECT 181.825 0.52 182.085 2.485 ;
      RECT 182.11 190.585 182.31 191.315 ;
      RECT 183.355 0.17 184.125 0.43 ;
      RECT 183.865 0.17 184.125 10.48 ;
      RECT 183.355 0.17 183.615 10.99 ;
      RECT 182.605 190.585 182.805 191.315 ;
      RECT 183.105 190.585 183.305 191.315 ;
      RECT 183.605 190.585 183.805 191.315 ;
      RECT 184.1 190.585 184.3 191.315 ;
      RECT 185.395 0.17 186.165 0.43 ;
      RECT 185.395 0.17 185.655 11.5 ;
      RECT 185.905 0.17 186.165 11.5 ;
      RECT 184.92 190.585 185.12 191.315 ;
      RECT 185.415 190.585 185.615 191.315 ;
      RECT 186.415 0.17 187.185 0.94 ;
      RECT 186.415 0.17 186.675 12.9 ;
      RECT 186.925 0.17 187.185 12.9 ;
      RECT 185.915 190.585 186.115 191.315 ;
      RECT 186.415 190.585 186.615 191.315 ;
      RECT 186.91 190.585 187.11 191.315 ;
      RECT 187.435 0.52 187.695 5.815 ;
      RECT 188.29 0.52 188.55 5.16 ;
      RECT 188.29 4.9 189.07 5.16 ;
      RECT 188.81 4.9 189.07 6.64 ;
      RECT 187.73 190.585 187.93 191.315 ;
      RECT 188.225 190.585 188.425 191.315 ;
      RECT 188.725 190.585 188.925 191.315 ;
      RECT 189.225 190.585 189.425 191.315 ;
      RECT 189.72 190.585 189.92 191.315 ;
      RECT 190.54 190.585 190.74 191.315 ;
      RECT 191.035 190.585 191.235 191.315 ;
      RECT 191.535 190.585 191.735 191.315 ;
      RECT 191.69 0.52 191.95 2.335 ;
      RECT 192.035 190.585 192.235 191.315 ;
      RECT 192.2 0.52 192.46 14.11 ;
      RECT 192.53 190.585 192.73 191.315 ;
      RECT 193.575 0.17 194.345 0.94 ;
      RECT 194.085 0.17 194.345 8.7 ;
      RECT 193.575 0.17 193.835 12.9 ;
      RECT 193.065 0.52 193.325 2.485 ;
      RECT 193.35 190.585 193.55 191.315 ;
      RECT 194.595 0.17 195.365 0.43 ;
      RECT 195.105 0.17 195.365 10.48 ;
      RECT 194.595 0.17 194.855 10.99 ;
      RECT 193.845 190.585 194.045 191.315 ;
      RECT 194.345 190.585 194.545 191.315 ;
      RECT 194.845 190.585 195.045 191.315 ;
      RECT 195.34 190.585 195.54 191.315 ;
      RECT 196.635 0.17 197.405 0.43 ;
      RECT 196.635 0.17 196.895 11.5 ;
      RECT 197.145 0.17 197.405 11.5 ;
      RECT 196.16 190.585 196.36 191.315 ;
      RECT 196.655 190.585 196.855 191.315 ;
      RECT 197.655 0.17 198.425 0.94 ;
      RECT 197.655 0.17 197.915 12.9 ;
      RECT 198.165 0.17 198.425 12.9 ;
      RECT 197.155 190.585 197.355 191.315 ;
      RECT 197.655 190.585 197.855 191.315 ;
      RECT 198.15 190.585 198.35 191.315 ;
      RECT 198.675 0.52 198.935 5.815 ;
      RECT 199.53 0.52 199.79 5.16 ;
      RECT 199.53 4.9 200.31 5.16 ;
      RECT 200.05 4.9 200.31 6.64 ;
      RECT 198.97 190.585 199.17 191.315 ;
      RECT 199.465 190.585 199.665 191.315 ;
      RECT 199.965 190.585 200.165 191.315 ;
      RECT 200.465 190.585 200.665 191.315 ;
      RECT 200.96 190.585 201.16 191.315 ;
      RECT 201.78 190.585 201.98 191.315 ;
      RECT 202.275 190.585 202.475 191.315 ;
      RECT 202.775 190.585 202.975 191.315 ;
      RECT 202.93 0.52 203.19 2.335 ;
      RECT 203.275 190.585 203.475 191.315 ;
      RECT 203.44 0.52 203.7 14.11 ;
      RECT 203.77 190.585 203.97 191.315 ;
      RECT 204.815 0.17 205.585 0.94 ;
      RECT 205.325 0.17 205.585 8.7 ;
      RECT 204.815 0.17 205.075 12.9 ;
      RECT 204.305 0.52 204.565 2.485 ;
      RECT 204.59 190.585 204.79 191.315 ;
      RECT 205.835 0.17 206.605 0.43 ;
      RECT 206.345 0.17 206.605 10.48 ;
      RECT 205.835 0.17 206.095 10.99 ;
      RECT 205.085 190.585 205.285 191.315 ;
      RECT 205.585 190.585 205.785 191.315 ;
      RECT 206.085 190.585 206.285 191.315 ;
      RECT 206.58 190.585 206.78 191.315 ;
      RECT 207.875 0.17 208.645 0.43 ;
      RECT 207.875 0.17 208.135 11.5 ;
      RECT 208.385 0.17 208.645 11.5 ;
      RECT 207.4 190.585 207.6 191.315 ;
      RECT 207.895 190.585 208.095 191.315 ;
      RECT 208.895 0.17 209.665 0.94 ;
      RECT 208.895 0.17 209.155 12.9 ;
      RECT 209.405 0.17 209.665 12.9 ;
      RECT 208.395 190.585 208.595 191.315 ;
      RECT 208.895 190.585 209.095 191.315 ;
      RECT 209.39 190.585 209.59 191.315 ;
      RECT 209.915 0.52 210.175 5.815 ;
      RECT 210.77 0.52 211.03 5.16 ;
      RECT 210.77 4.9 211.55 5.16 ;
      RECT 211.29 4.9 211.55 6.64 ;
      RECT 210.21 190.585 210.41 191.315 ;
      RECT 210.705 190.585 210.905 191.315 ;
      RECT 211.205 190.585 211.405 191.315 ;
      RECT 211.705 190.585 211.905 191.315 ;
      RECT 212.2 190.585 212.4 191.315 ;
      RECT 213.02 190.585 213.22 191.315 ;
      RECT 213.515 190.585 213.715 191.315 ;
      RECT 214.015 190.585 214.215 191.315 ;
      RECT 214.17 0.52 214.43 2.335 ;
      RECT 214.515 190.585 214.715 191.315 ;
      RECT 214.68 0.52 214.94 14.11 ;
      RECT 215.01 190.585 215.21 191.315 ;
      RECT 216.055 0.17 216.825 0.94 ;
      RECT 216.565 0.17 216.825 8.7 ;
      RECT 216.055 0.17 216.315 12.9 ;
      RECT 215.545 0.52 215.805 2.485 ;
      RECT 215.83 190.585 216.03 191.315 ;
      RECT 217.075 0.17 217.845 0.43 ;
      RECT 217.585 0.17 217.845 10.48 ;
      RECT 217.075 0.17 217.335 10.99 ;
      RECT 216.325 190.585 216.525 191.315 ;
      RECT 216.825 190.585 217.025 191.315 ;
      RECT 217.325 190.585 217.525 191.315 ;
      RECT 217.82 190.585 218.02 191.315 ;
      RECT 219.115 0.17 219.885 0.43 ;
      RECT 219.115 0.17 219.375 11.5 ;
      RECT 219.625 0.17 219.885 11.5 ;
      RECT 218.64 190.585 218.84 191.315 ;
      RECT 219.135 190.585 219.335 191.315 ;
      RECT 220.135 0.17 220.905 0.94 ;
      RECT 220.135 0.17 220.395 12.9 ;
      RECT 220.645 0.17 220.905 12.9 ;
      RECT 219.635 190.585 219.835 191.315 ;
      RECT 220.135 190.585 220.335 191.315 ;
      RECT 220.63 190.585 220.83 191.315 ;
      RECT 221.155 0.52 221.415 5.815 ;
      RECT 222.01 0.52 222.27 5.16 ;
      RECT 222.01 4.9 222.79 5.16 ;
      RECT 222.53 4.9 222.79 6.64 ;
      RECT 221.45 190.585 221.65 191.315 ;
      RECT 221.945 190.585 222.145 191.315 ;
      RECT 222.445 190.585 222.645 191.315 ;
      RECT 222.945 190.585 223.145 191.315 ;
      RECT 223.44 190.585 223.64 191.315 ;
      RECT 224.26 190.585 224.46 191.315 ;
      RECT 224.755 190.585 224.955 191.315 ;
      RECT 225.255 190.585 225.455 191.315 ;
      RECT 225.41 0.52 225.67 2.335 ;
      RECT 225.755 190.585 225.955 191.315 ;
      RECT 225.92 0.52 226.18 14.11 ;
      RECT 226.25 190.585 226.45 191.315 ;
      RECT 227.295 0.17 228.065 0.94 ;
      RECT 227.805 0.17 228.065 8.7 ;
      RECT 227.295 0.17 227.555 12.9 ;
      RECT 226.785 0.52 227.045 2.485 ;
      RECT 227.07 190.585 227.27 191.315 ;
      RECT 228.315 0.17 229.085 0.43 ;
      RECT 228.825 0.17 229.085 10.48 ;
      RECT 228.315 0.17 228.575 10.99 ;
      RECT 227.565 190.585 227.765 191.315 ;
      RECT 228.065 190.585 228.265 191.315 ;
      RECT 228.565 190.585 228.765 191.315 ;
      RECT 229.06 190.585 229.26 191.315 ;
      RECT 230.355 0.17 231.125 0.43 ;
      RECT 230.355 0.17 230.615 11.5 ;
      RECT 230.865 0.17 231.125 11.5 ;
      RECT 229.88 190.585 230.08 191.315 ;
      RECT 230.375 190.585 230.575 191.315 ;
      RECT 231.375 0.17 232.145 0.94 ;
      RECT 231.375 0.17 231.635 12.9 ;
      RECT 231.885 0.17 232.145 12.9 ;
      RECT 230.875 190.585 231.075 191.315 ;
      RECT 231.375 190.585 231.575 191.315 ;
      RECT 231.87 190.585 232.07 191.315 ;
      RECT 232.395 0.52 232.655 5.815 ;
      RECT 233.25 0.52 233.51 5.16 ;
      RECT 233.25 4.9 234.03 5.16 ;
      RECT 233.77 4.9 234.03 6.64 ;
      RECT 232.69 190.585 232.89 191.315 ;
      RECT 233.185 190.585 233.385 191.315 ;
      RECT 233.685 190.585 233.885 191.315 ;
      RECT 234.185 190.585 234.385 191.315 ;
      RECT 234.68 190.585 234.88 191.315 ;
      RECT 235.5 190.585 235.7 191.315 ;
      RECT 236.495 45.465 236.695 191.315 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 113.59 0 113.83 191.34 ;
      RECT 116.65 0 116.89 191.34 ;
      RECT 118.18 0 118.42 191.34 ;
      RECT 125.31 0 132.19 191.34 ;
      RECT 133.48 0 134.23 191.34 ;
      RECT 0 0 3.03 191.34 ;
      RECT 4.655 0.17 9.505 191.34 ;
      RECT 11.65 0 14.27 191.34 ;
      RECT 15.895 0.17 20.745 191.34 ;
      RECT 22.89 0 25.51 191.34 ;
      RECT 27.135 0.17 31.985 191.34 ;
      RECT 34.13 0 36.75 191.34 ;
      RECT 38.375 0.17 43.225 191.34 ;
      RECT 45.37 0 47.99 191.34 ;
      RECT 49.615 0.17 54.465 191.34 ;
      RECT 56.61 0 59.23 191.34 ;
      RECT 60.855 0.17 65.705 191.34 ;
      RECT 67.85 0 70.47 191.34 ;
      RECT 72.095 0.17 76.945 191.34 ;
      RECT 79.09 0 81.71 191.34 ;
      RECT 83.335 0.17 88.185 191.34 ;
      RECT 90.33 0 102.11 191.34 ;
      RECT 104.4 0.17 110.78 191.34 ;
      RECT 112.05 0.3 112.31 191.34 ;
      RECT 113.58 0.3 113.84 191.34 ;
      RECT 116.64 0.3 116.9 191.34 ;
      RECT 118.17 0.3 118.43 191.34 ;
      RECT 119.71 0.17 120.98 191.34 ;
      RECT 119.7 0.3 120.98 191.34 ;
      RECT 125.31 0.3 132.2 191.34 ;
      RECT 133.47 0.3 134.24 191.34 ;
      RECT 135.01 0 146.47 191.34 ;
      RECT 135 0.17 146.47 191.34 ;
      RECT 148.615 0.17 153.465 191.34 ;
      RECT 155.09 0 157.71 191.34 ;
      RECT 159.855 0.17 164.705 191.34 ;
      RECT 166.33 0 168.95 191.34 ;
      RECT 171.095 0.17 175.945 191.34 ;
      RECT 177.57 0 180.19 191.34 ;
      RECT 182.335 0.17 187.185 191.34 ;
      RECT 188.81 0 191.43 191.34 ;
      RECT 193.575 0.17 198.425 191.34 ;
      RECT 200.05 0 202.67 191.34 ;
      RECT 204.815 0.17 209.665 191.34 ;
      RECT 211.29 0 213.91 191.34 ;
      RECT 216.055 0.17 220.905 191.34 ;
      RECT 222.53 0 225.15 191.34 ;
      RECT 227.295 0.17 232.145 191.34 ;
      RECT 233.77 0 236.8 191.34 ;
      RECT 0 0.52 236.8 191.34 ;
      RECT 4.665 0 9.495 191.34 ;
      RECT 15.905 0 20.735 191.34 ;
      RECT 27.145 0 31.975 191.34 ;
      RECT 38.385 0 43.215 191.34 ;
      RECT 49.625 0 54.455 191.34 ;
      RECT 60.865 0 65.695 191.34 ;
      RECT 72.105 0 76.935 191.34 ;
      RECT 83.345 0 88.175 191.34 ;
      RECT 104.4 0 110.77 191.34 ;
      RECT 119.71 0 120.97 191.34 ;
      RECT 148.625 0 153.455 191.34 ;
      RECT 159.865 0 164.695 191.34 ;
      RECT 171.105 0 175.935 191.34 ;
      RECT 182.345 0 187.175 191.34 ;
      RECT 193.585 0 198.415 191.34 ;
      RECT 204.825 0 209.655 191.34 ;
      RECT 216.065 0 220.895 191.34 ;
      RECT 227.305 0 232.135 191.34 ;
      RECT 112.06 0 112.3 191.34 ;
    LAYER Metal3 ;
      RECT 0 0 236.8 191.34 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 39.085 9.62 45.205 ;
      RECT 0 0 4 191.34 ;
      RECT 7.33 0 9.62 191.34 ;
      RECT 12.95 39.085 20.86 45.205 ;
      RECT 12.95 0 15.24 191.34 ;
      RECT 18.57 0 20.86 191.34 ;
      RECT 24.19 39.085 32.1 45.205 ;
      RECT 24.19 0 26.48 191.34 ;
      RECT 29.81 0 32.1 191.34 ;
      RECT 35.43 39.085 43.34 45.205 ;
      RECT 35.43 0 37.72 191.34 ;
      RECT 41.05 0 43.34 191.34 ;
      RECT 46.67 39.085 54.58 45.205 ;
      RECT 46.67 0 48.96 191.34 ;
      RECT 52.29 0 54.58 191.34 ;
      RECT 57.91 39.085 65.82 45.205 ;
      RECT 57.91 0 60.2 191.34 ;
      RECT 63.53 0 65.82 191.34 ;
      RECT 69.15 39.085 77.06 45.205 ;
      RECT 69.15 0 71.44 191.34 ;
      RECT 74.77 0 77.06 191.34 ;
      RECT 80.39 39.085 88.3 45.205 ;
      RECT 80.39 0 82.68 191.34 ;
      RECT 86.01 0 88.3 191.34 ;
      RECT 91.63 0 98.71 191.34 ;
      RECT 102.04 0 103.86 191.34 ;
      RECT 107.19 0 109.01 191.34 ;
      RECT 112.34 0 114.16 191.34 ;
      RECT 117.49 0 119.31 191.34 ;
      RECT 122.64 0 124.46 191.34 ;
      RECT 148.5 39.085 156.41 45.205 ;
      RECT 148.5 0 150.79 191.34 ;
      RECT 154.12 0 156.41 191.34 ;
      RECT 159.74 39.085 167.65 45.205 ;
      RECT 159.74 0 162.03 191.34 ;
      RECT 165.36 0 167.65 191.34 ;
      RECT 170.98 39.085 178.89 45.205 ;
      RECT 170.98 0 173.27 191.34 ;
      RECT 176.6 0 178.89 191.34 ;
      RECT 182.22 39.085 190.13 45.205 ;
      RECT 182.22 0 184.51 191.34 ;
      RECT 187.84 0 190.13 191.34 ;
      RECT 193.46 39.085 201.37 45.205 ;
      RECT 193.46 0 195.75 191.34 ;
      RECT 199.08 0 201.37 191.34 ;
      RECT 204.7 39.085 212.61 45.205 ;
      RECT 204.7 0 206.99 191.34 ;
      RECT 210.32 0 212.61 191.34 ;
      RECT 215.94 39.085 223.85 45.205 ;
      RECT 215.94 0 218.23 191.34 ;
      RECT 221.56 0 223.85 191.34 ;
      RECT 227.18 39.085 236.8 45.205 ;
      RECT 227.18 0 229.47 191.34 ;
      RECT 232.8 0 236.8 191.34 ;
      RECT 127.79 0 129.61 191.34 ;
      RECT 132.94 0 134.76 191.34 ;
      RECT 138.09 0 145.17 191.34 ;
  END
END RM_IHPSG13_1P_512x16_c2_bm_bist

END LIBRARY
