# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Thu Aug 21 20:48:28 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_1024x32_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_1024x32_c2_bm_bist 0 0 ;
  SIZE 416.64 BY 336.46 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 244.49 0 244.75 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171.89 0 172.15 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 243.635 0 243.895 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.745 0 173.005 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 236.65 0 236.91 0.26 ;
    END
  END A_BM[16]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.73 0 179.99 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 238.025 0 238.285 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.355 0 178.615 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 237.16 0 237.42 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.22 0 179.48 0.26 ;
    END
  END A_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 403.95 0 406.76 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.71 0 395.52 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 381.47 0 384.28 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.23 0 373.04 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.99 0 361.8 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.75 0 350.56 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 336.51 0 339.32 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.27 0 328.08 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.03 0 316.84 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.79 0 305.6 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 291.55 0 294.36 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.31 0 283.12 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.07 0 271.88 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 257.83 0 260.64 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.59 0 249.4 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.35 0 238.16 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.94 0 227.75 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.64 0 217.45 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 199.19 0 202 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 188.89 0 191.7 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.48 0 181.29 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.24 0 170.05 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156 0 158.81 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 144.76 0 147.57 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.52 0 136.33 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.28 0 125.09 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.04 0 113.85 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.8 0 102.61 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 336.46 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 0 412.38 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 0 401.14 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 0 389.9 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 0 378.66 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 0 367.42 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 0 356.18 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 0 344.94 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 0 333.7 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 0 322.46 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 0 311.22 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 0 299.98 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 0 288.74 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 0 277.5 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 0 266.26 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 0 255.02 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 0 243.78 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.79 0 222.6 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.49 0 212.3 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 204.34 0 207.15 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 194.04 0 196.85 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 0 175.67 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 0 164.43 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 0 153.19 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 0 141.95 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 0 130.71 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 0 119.47 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 0 108.23 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 0 96.99 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 38.825 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 45.465 412.38 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 45.465 401.14 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 45.465 389.9 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 45.465 378.66 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 45.465 367.42 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 45.465 356.18 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 45.465 344.94 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 45.465 333.7 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 45.465 322.46 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 45.465 311.22 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 45.465 299.98 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 45.465 288.74 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 45.465 277.5 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 45.465 266.26 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 45.465 255.02 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 45.465 243.78 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 45.465 175.67 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 45.465 164.43 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 45.465 153.19 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 45.465 141.95 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 45.465 130.71 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 45.465 119.47 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 45.465 108.23 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 45.465 96.99 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 45.465 85.75 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 45.465 74.51 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 45.465 63.27 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 45.465 52.03 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 45.465 40.79 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 45.465 29.55 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 45.465 18.31 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 45.465 7.07 336.46 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 255.73 0 255.99 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.65 0 160.91 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 254.875 0 255.135 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.505 0 161.765 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 247.89 0 248.15 0.26 ;
    END
  END A_BM[17]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.49 0 168.75 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.265 0 249.525 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.115 0 167.375 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.4 0 248.66 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.98 0 168.24 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.97 0 267.23 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 149.41 0 149.67 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.115 0 266.375 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.265 0 150.525 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.13 0 259.39 0.26 ;
    END
  END A_BM[18]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.25 0 157.51 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 260.505 0 260.765 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.875 0 156.135 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.64 0 259.9 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.74 0 157 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 278.21 0 278.47 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 138.17 0 138.43 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.355 0 277.615 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 139.025 0 139.285 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 270.37 0 270.63 0.26 ;
    END
  END A_BM[19]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.01 0 146.27 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 271.745 0 272.005 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.635 0 144.895 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 270.88 0 271.14 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.5 0 145.76 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 289.45 0 289.71 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.93 0 127.19 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 288.595 0 288.855 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 127.785 0 128.045 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 281.61 0 281.87 0.26 ;
    END
  END A_BM[20]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.77 0 135.03 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.985 0 283.245 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.395 0 133.655 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.12 0 282.38 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.26 0 134.52 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 300.69 0 300.95 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.69 0 115.95 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 299.835 0 300.095 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.545 0 116.805 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 292.85 0 293.11 0.26 ;
    END
  END A_BM[21]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.53 0 123.79 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.225 0 294.485 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.155 0 122.415 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.36 0 293.62 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.02 0 123.28 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.93 0 312.19 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.45 0 104.71 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.075 0 311.335 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 105.305 0 105.565 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.09 0 304.35 0.26 ;
    END
  END A_BM[22]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.29 0 112.55 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 305.465 0 305.725 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.915 0 111.175 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.6 0 304.86 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.78 0 112.04 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 323.17 0 323.43 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 93.21 0 93.47 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 322.315 0 322.575 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 94.065 0 94.325 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.33 0 315.59 0.26 ;
    END
  END A_BM[23]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.05 0 101.31 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 316.705 0 316.965 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.675 0 99.935 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.84 0 316.1 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.54 0 100.8 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.41 0 334.67 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.97 0 82.23 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.555 0 333.815 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.825 0 83.085 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 326.57 0 326.83 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.81 0 90.07 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.945 0 328.205 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.435 0 88.695 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.08 0 327.34 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.3 0 89.56 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 345.65 0 345.91 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.73 0 70.99 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 344.795 0 345.055 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 71.585 0 71.845 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.81 0 338.07 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.57 0 78.83 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.185 0 339.445 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.195 0 77.455 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.32 0 338.58 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.06 0 78.32 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.89 0 357.15 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 59.49 0 59.75 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.035 0 356.295 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.345 0 60.605 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.05 0 349.31 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.33 0 67.59 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 350.425 0 350.685 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 65.955 0 66.215 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.56 0 349.82 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.82 0 67.08 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.13 0 368.39 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 48.25 0 48.51 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 367.275 0 367.535 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 49.105 0 49.365 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.29 0 360.55 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.09 0 56.35 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 361.665 0 361.925 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.715 0 54.975 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.8 0 361.06 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.58 0 55.84 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.37 0 379.63 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.01 0 37.27 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.515 0 378.775 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.865 0 38.125 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.53 0 371.79 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.85 0 45.11 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.905 0 373.165 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 43.475 0 43.735 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.04 0 372.3 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.34 0 44.6 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.61 0 390.87 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 25.77 0 26.03 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 389.755 0 390.015 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 26.625 0 26.885 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.77 0 383.03 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.61 0 33.87 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.145 0 384.405 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.235 0 32.495 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 383.28 0 383.54 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.1 0 33.36 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.85 0 402.11 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.53 0 14.79 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.995 0 401.255 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.385 0 15.645 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.01 0 394.27 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.37 0 22.63 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 395.385 0 395.645 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.995 0 21.255 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.52 0 394.78 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 21.86 0 22.12 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 413.09 0 413.35 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.29 0 3.55 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 412.235 0 412.495 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.145 0 4.405 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.25 0 405.51 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.13 0 11.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 406.625 0 406.885 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.755 0 10.015 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.76 0 406.02 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.62 0 10.88 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 45.223301 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.52 0 204.78 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.184466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 209.11 0 209.37 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 39.656958 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.01 0 204.27 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.618123 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 208.6 0 208.86 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.17 0 212.43 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.68 0 212.94 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.15 0 211.41 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.66 0 211.92 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.63754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.72 0 214.98 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.317152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.21 0 214.47 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 70.245955 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.7 0 213.96 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 68.925566 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.19 0 213.45 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 55.436893 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.28 0 192.54 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 54.065721 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.79 0 193.05 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 62.724919 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.3 0 193.56 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.404531 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.81 0 194.07 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.740105 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 222.37 0 222.63 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.204381 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 222.88 0 223.14 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2633 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.963157 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.27 0 217.53 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0083 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.693552 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.78 0 218.04 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.48 0 202.74 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.796863 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.05 0 206.31 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.54 0 205.8 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.99 0 203.25 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 18.532819 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.41 0 224.67 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 203.31695 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.885 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.213636 LAYER Metal2 ;
      ANTENNAMAXAREACAR 17.563993 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.03 0 205.29 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.95 0 201.21 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.58 0 207.84 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.07 0 207.33 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 201.46 0 201.72 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 416.64 336.46 ;
    LAYER Metal2 ;
      RECT 0.105 45.465 0.305 336.435 ;
      RECT 1.1 335.705 1.3 336.435 ;
      RECT 3.29 0.52 3.55 5.16 ;
      RECT 2.77 4.9 3.55 5.16 ;
      RECT 2.77 4.9 3.03 6.64 ;
      RECT 1.92 335.705 2.12 336.435 ;
      RECT 2.415 335.705 2.615 336.435 ;
      RECT 2.915 335.705 3.115 336.435 ;
      RECT 3.415 335.705 3.615 336.435 ;
      RECT 3.91 335.705 4.11 336.435 ;
      RECT 4.655 0.17 5.425 0.94 ;
      RECT 4.655 0.17 4.915 12.9 ;
      RECT 5.165 0.17 5.425 12.9 ;
      RECT 4.145 0.52 4.405 5.815 ;
      RECT 4.73 335.705 4.93 336.435 ;
      RECT 5.675 0.17 6.445 0.43 ;
      RECT 5.675 0.17 5.935 11.5 ;
      RECT 6.185 0.17 6.445 11.5 ;
      RECT 5.225 335.705 5.425 336.435 ;
      RECT 5.725 335.705 5.925 336.435 ;
      RECT 6.225 335.705 6.425 336.435 ;
      RECT 7.715 0.17 8.485 0.43 ;
      RECT 7.715 0.17 7.975 10.48 ;
      RECT 8.225 0.17 8.485 10.99 ;
      RECT 6.72 335.705 6.92 336.435 ;
      RECT 7.54 335.705 7.74 336.435 ;
      RECT 8.735 0.17 9.505 0.94 ;
      RECT 8.735 0.17 8.995 8.7 ;
      RECT 9.245 0.17 9.505 12.9 ;
      RECT 8.035 335.705 8.235 336.435 ;
      RECT 8.535 335.705 8.735 336.435 ;
      RECT 9.035 335.705 9.235 336.435 ;
      RECT 9.53 335.705 9.73 336.435 ;
      RECT 9.755 0.52 10.015 2.485 ;
      RECT 10.35 335.705 10.55 336.435 ;
      RECT 10.62 0.52 10.88 14.11 ;
      RECT 10.845 335.705 11.045 336.435 ;
      RECT 11.13 0.52 11.39 2.335 ;
      RECT 11.345 335.705 11.545 336.435 ;
      RECT 11.845 335.705 12.045 336.435 ;
      RECT 12.34 335.705 12.54 336.435 ;
      RECT 14.53 0.52 14.79 5.16 ;
      RECT 14.01 4.9 14.79 5.16 ;
      RECT 14.01 4.9 14.27 6.64 ;
      RECT 13.16 335.705 13.36 336.435 ;
      RECT 13.655 335.705 13.855 336.435 ;
      RECT 14.155 335.705 14.355 336.435 ;
      RECT 14.655 335.705 14.855 336.435 ;
      RECT 15.15 335.705 15.35 336.435 ;
      RECT 15.895 0.17 16.665 0.94 ;
      RECT 15.895 0.17 16.155 12.9 ;
      RECT 16.405 0.17 16.665 12.9 ;
      RECT 15.385 0.52 15.645 5.815 ;
      RECT 15.97 335.705 16.17 336.435 ;
      RECT 16.915 0.17 17.685 0.43 ;
      RECT 16.915 0.17 17.175 11.5 ;
      RECT 17.425 0.17 17.685 11.5 ;
      RECT 16.465 335.705 16.665 336.435 ;
      RECT 16.965 335.705 17.165 336.435 ;
      RECT 17.465 335.705 17.665 336.435 ;
      RECT 18.955 0.17 19.725 0.43 ;
      RECT 18.955 0.17 19.215 10.48 ;
      RECT 19.465 0.17 19.725 10.99 ;
      RECT 17.96 335.705 18.16 336.435 ;
      RECT 18.78 335.705 18.98 336.435 ;
      RECT 19.975 0.17 20.745 0.94 ;
      RECT 19.975 0.17 20.235 8.7 ;
      RECT 20.485 0.17 20.745 12.9 ;
      RECT 19.275 335.705 19.475 336.435 ;
      RECT 19.775 335.705 19.975 336.435 ;
      RECT 20.275 335.705 20.475 336.435 ;
      RECT 20.77 335.705 20.97 336.435 ;
      RECT 20.995 0.52 21.255 2.485 ;
      RECT 21.59 335.705 21.79 336.435 ;
      RECT 21.86 0.52 22.12 14.11 ;
      RECT 22.085 335.705 22.285 336.435 ;
      RECT 22.37 0.52 22.63 2.335 ;
      RECT 22.585 335.705 22.785 336.435 ;
      RECT 23.085 335.705 23.285 336.435 ;
      RECT 23.58 335.705 23.78 336.435 ;
      RECT 25.77 0.52 26.03 5.16 ;
      RECT 25.25 4.9 26.03 5.16 ;
      RECT 25.25 4.9 25.51 6.64 ;
      RECT 24.4 335.705 24.6 336.435 ;
      RECT 24.895 335.705 25.095 336.435 ;
      RECT 25.395 335.705 25.595 336.435 ;
      RECT 25.895 335.705 26.095 336.435 ;
      RECT 26.39 335.705 26.59 336.435 ;
      RECT 27.135 0.17 27.905 0.94 ;
      RECT 27.135 0.17 27.395 12.9 ;
      RECT 27.645 0.17 27.905 12.9 ;
      RECT 26.625 0.52 26.885 5.815 ;
      RECT 27.21 335.705 27.41 336.435 ;
      RECT 28.155 0.17 28.925 0.43 ;
      RECT 28.155 0.17 28.415 11.5 ;
      RECT 28.665 0.17 28.925 11.5 ;
      RECT 27.705 335.705 27.905 336.435 ;
      RECT 28.205 335.705 28.405 336.435 ;
      RECT 28.705 335.705 28.905 336.435 ;
      RECT 30.195 0.17 30.965 0.43 ;
      RECT 30.195 0.17 30.455 10.48 ;
      RECT 30.705 0.17 30.965 10.99 ;
      RECT 29.2 335.705 29.4 336.435 ;
      RECT 30.02 335.705 30.22 336.435 ;
      RECT 31.215 0.17 31.985 0.94 ;
      RECT 31.215 0.17 31.475 8.7 ;
      RECT 31.725 0.17 31.985 12.9 ;
      RECT 30.515 335.705 30.715 336.435 ;
      RECT 31.015 335.705 31.215 336.435 ;
      RECT 31.515 335.705 31.715 336.435 ;
      RECT 32.01 335.705 32.21 336.435 ;
      RECT 32.235 0.52 32.495 2.485 ;
      RECT 32.83 335.705 33.03 336.435 ;
      RECT 33.1 0.52 33.36 14.11 ;
      RECT 33.325 335.705 33.525 336.435 ;
      RECT 33.61 0.52 33.87 2.335 ;
      RECT 33.825 335.705 34.025 336.435 ;
      RECT 34.325 335.705 34.525 336.435 ;
      RECT 34.82 335.705 35.02 336.435 ;
      RECT 37.01 0.52 37.27 5.16 ;
      RECT 36.49 4.9 37.27 5.16 ;
      RECT 36.49 4.9 36.75 6.64 ;
      RECT 35.64 335.705 35.84 336.435 ;
      RECT 36.135 335.705 36.335 336.435 ;
      RECT 36.635 335.705 36.835 336.435 ;
      RECT 37.135 335.705 37.335 336.435 ;
      RECT 37.63 335.705 37.83 336.435 ;
      RECT 38.375 0.17 39.145 0.94 ;
      RECT 38.375 0.17 38.635 12.9 ;
      RECT 38.885 0.17 39.145 12.9 ;
      RECT 37.865 0.52 38.125 5.815 ;
      RECT 38.45 335.705 38.65 336.435 ;
      RECT 39.395 0.17 40.165 0.43 ;
      RECT 39.395 0.17 39.655 11.5 ;
      RECT 39.905 0.17 40.165 11.5 ;
      RECT 38.945 335.705 39.145 336.435 ;
      RECT 39.445 335.705 39.645 336.435 ;
      RECT 39.945 335.705 40.145 336.435 ;
      RECT 41.435 0.17 42.205 0.43 ;
      RECT 41.435 0.17 41.695 10.48 ;
      RECT 41.945 0.17 42.205 10.99 ;
      RECT 40.44 335.705 40.64 336.435 ;
      RECT 41.26 335.705 41.46 336.435 ;
      RECT 42.455 0.17 43.225 0.94 ;
      RECT 42.455 0.17 42.715 8.7 ;
      RECT 42.965 0.17 43.225 12.9 ;
      RECT 41.755 335.705 41.955 336.435 ;
      RECT 42.255 335.705 42.455 336.435 ;
      RECT 42.755 335.705 42.955 336.435 ;
      RECT 43.25 335.705 43.45 336.435 ;
      RECT 43.475 0.52 43.735 2.485 ;
      RECT 44.07 335.705 44.27 336.435 ;
      RECT 44.34 0.52 44.6 14.11 ;
      RECT 44.565 335.705 44.765 336.435 ;
      RECT 44.85 0.52 45.11 2.335 ;
      RECT 45.065 335.705 45.265 336.435 ;
      RECT 45.565 335.705 45.765 336.435 ;
      RECT 46.06 335.705 46.26 336.435 ;
      RECT 48.25 0.52 48.51 5.16 ;
      RECT 47.73 4.9 48.51 5.16 ;
      RECT 47.73 4.9 47.99 6.64 ;
      RECT 46.88 335.705 47.08 336.435 ;
      RECT 47.375 335.705 47.575 336.435 ;
      RECT 47.875 335.705 48.075 336.435 ;
      RECT 48.375 335.705 48.575 336.435 ;
      RECT 48.87 335.705 49.07 336.435 ;
      RECT 49.615 0.17 50.385 0.94 ;
      RECT 49.615 0.17 49.875 12.9 ;
      RECT 50.125 0.17 50.385 12.9 ;
      RECT 49.105 0.52 49.365 5.815 ;
      RECT 49.69 335.705 49.89 336.435 ;
      RECT 50.635 0.17 51.405 0.43 ;
      RECT 50.635 0.17 50.895 11.5 ;
      RECT 51.145 0.17 51.405 11.5 ;
      RECT 50.185 335.705 50.385 336.435 ;
      RECT 50.685 335.705 50.885 336.435 ;
      RECT 51.185 335.705 51.385 336.435 ;
      RECT 52.675 0.17 53.445 0.43 ;
      RECT 52.675 0.17 52.935 10.48 ;
      RECT 53.185 0.17 53.445 10.99 ;
      RECT 51.68 335.705 51.88 336.435 ;
      RECT 52.5 335.705 52.7 336.435 ;
      RECT 53.695 0.17 54.465 0.94 ;
      RECT 53.695 0.17 53.955 8.7 ;
      RECT 54.205 0.17 54.465 12.9 ;
      RECT 52.995 335.705 53.195 336.435 ;
      RECT 53.495 335.705 53.695 336.435 ;
      RECT 53.995 335.705 54.195 336.435 ;
      RECT 54.49 335.705 54.69 336.435 ;
      RECT 54.715 0.52 54.975 2.485 ;
      RECT 55.31 335.705 55.51 336.435 ;
      RECT 55.58 0.52 55.84 14.11 ;
      RECT 55.805 335.705 56.005 336.435 ;
      RECT 56.09 0.52 56.35 2.335 ;
      RECT 56.305 335.705 56.505 336.435 ;
      RECT 56.805 335.705 57.005 336.435 ;
      RECT 57.3 335.705 57.5 336.435 ;
      RECT 59.49 0.52 59.75 5.16 ;
      RECT 58.97 4.9 59.75 5.16 ;
      RECT 58.97 4.9 59.23 6.64 ;
      RECT 58.12 335.705 58.32 336.435 ;
      RECT 58.615 335.705 58.815 336.435 ;
      RECT 59.115 335.705 59.315 336.435 ;
      RECT 59.615 335.705 59.815 336.435 ;
      RECT 60.11 335.705 60.31 336.435 ;
      RECT 60.855 0.17 61.625 0.94 ;
      RECT 60.855 0.17 61.115 12.9 ;
      RECT 61.365 0.17 61.625 12.9 ;
      RECT 60.345 0.52 60.605 5.815 ;
      RECT 60.93 335.705 61.13 336.435 ;
      RECT 61.875 0.17 62.645 0.43 ;
      RECT 61.875 0.17 62.135 11.5 ;
      RECT 62.385 0.17 62.645 11.5 ;
      RECT 61.425 335.705 61.625 336.435 ;
      RECT 61.925 335.705 62.125 336.435 ;
      RECT 62.425 335.705 62.625 336.435 ;
      RECT 63.915 0.17 64.685 0.43 ;
      RECT 63.915 0.17 64.175 10.48 ;
      RECT 64.425 0.17 64.685 10.99 ;
      RECT 62.92 335.705 63.12 336.435 ;
      RECT 63.74 335.705 63.94 336.435 ;
      RECT 64.935 0.17 65.705 0.94 ;
      RECT 64.935 0.17 65.195 8.7 ;
      RECT 65.445 0.17 65.705 12.9 ;
      RECT 64.235 335.705 64.435 336.435 ;
      RECT 64.735 335.705 64.935 336.435 ;
      RECT 65.235 335.705 65.435 336.435 ;
      RECT 65.73 335.705 65.93 336.435 ;
      RECT 65.955 0.52 66.215 2.485 ;
      RECT 66.55 335.705 66.75 336.435 ;
      RECT 66.82 0.52 67.08 14.11 ;
      RECT 67.045 335.705 67.245 336.435 ;
      RECT 67.33 0.52 67.59 2.335 ;
      RECT 67.545 335.705 67.745 336.435 ;
      RECT 68.045 335.705 68.245 336.435 ;
      RECT 68.54 335.705 68.74 336.435 ;
      RECT 70.73 0.52 70.99 5.16 ;
      RECT 70.21 4.9 70.99 5.16 ;
      RECT 70.21 4.9 70.47 6.64 ;
      RECT 69.36 335.705 69.56 336.435 ;
      RECT 69.855 335.705 70.055 336.435 ;
      RECT 70.355 335.705 70.555 336.435 ;
      RECT 70.855 335.705 71.055 336.435 ;
      RECT 71.35 335.705 71.55 336.435 ;
      RECT 72.095 0.17 72.865 0.94 ;
      RECT 72.095 0.17 72.355 12.9 ;
      RECT 72.605 0.17 72.865 12.9 ;
      RECT 71.585 0.52 71.845 5.815 ;
      RECT 72.17 335.705 72.37 336.435 ;
      RECT 73.115 0.17 73.885 0.43 ;
      RECT 73.115 0.17 73.375 11.5 ;
      RECT 73.625 0.17 73.885 11.5 ;
      RECT 72.665 335.705 72.865 336.435 ;
      RECT 73.165 335.705 73.365 336.435 ;
      RECT 73.665 335.705 73.865 336.435 ;
      RECT 75.155 0.17 75.925 0.43 ;
      RECT 75.155 0.17 75.415 10.48 ;
      RECT 75.665 0.17 75.925 10.99 ;
      RECT 74.16 335.705 74.36 336.435 ;
      RECT 74.98 335.705 75.18 336.435 ;
      RECT 76.175 0.17 76.945 0.94 ;
      RECT 76.175 0.17 76.435 8.7 ;
      RECT 76.685 0.17 76.945 12.9 ;
      RECT 75.475 335.705 75.675 336.435 ;
      RECT 75.975 335.705 76.175 336.435 ;
      RECT 76.475 335.705 76.675 336.435 ;
      RECT 76.97 335.705 77.17 336.435 ;
      RECT 77.195 0.52 77.455 2.485 ;
      RECT 77.79 335.705 77.99 336.435 ;
      RECT 78.06 0.52 78.32 14.11 ;
      RECT 78.285 335.705 78.485 336.435 ;
      RECT 78.57 0.52 78.83 2.335 ;
      RECT 78.785 335.705 78.985 336.435 ;
      RECT 79.285 335.705 79.485 336.435 ;
      RECT 79.78 335.705 79.98 336.435 ;
      RECT 81.97 0.52 82.23 5.16 ;
      RECT 81.45 4.9 82.23 5.16 ;
      RECT 81.45 4.9 81.71 6.64 ;
      RECT 80.6 335.705 80.8 336.435 ;
      RECT 81.095 335.705 81.295 336.435 ;
      RECT 81.595 335.705 81.795 336.435 ;
      RECT 82.095 335.705 82.295 336.435 ;
      RECT 82.59 335.705 82.79 336.435 ;
      RECT 83.335 0.17 84.105 0.94 ;
      RECT 83.335 0.17 83.595 12.9 ;
      RECT 83.845 0.17 84.105 12.9 ;
      RECT 82.825 0.52 83.085 5.815 ;
      RECT 83.41 335.705 83.61 336.435 ;
      RECT 84.355 0.17 85.125 0.43 ;
      RECT 84.355 0.17 84.615 11.5 ;
      RECT 84.865 0.17 85.125 11.5 ;
      RECT 83.905 335.705 84.105 336.435 ;
      RECT 84.405 335.705 84.605 336.435 ;
      RECT 84.905 335.705 85.105 336.435 ;
      RECT 86.395 0.17 87.165 0.43 ;
      RECT 86.395 0.17 86.655 10.48 ;
      RECT 86.905 0.17 87.165 10.99 ;
      RECT 85.4 335.705 85.6 336.435 ;
      RECT 86.22 335.705 86.42 336.435 ;
      RECT 87.415 0.17 88.185 0.94 ;
      RECT 87.415 0.17 87.675 8.7 ;
      RECT 87.925 0.17 88.185 12.9 ;
      RECT 86.715 335.705 86.915 336.435 ;
      RECT 87.215 335.705 87.415 336.435 ;
      RECT 87.715 335.705 87.915 336.435 ;
      RECT 88.21 335.705 88.41 336.435 ;
      RECT 88.435 0.52 88.695 2.485 ;
      RECT 89.03 335.705 89.23 336.435 ;
      RECT 89.3 0.52 89.56 14.11 ;
      RECT 89.525 335.705 89.725 336.435 ;
      RECT 89.81 0.52 90.07 2.335 ;
      RECT 90.025 335.705 90.225 336.435 ;
      RECT 90.525 335.705 90.725 336.435 ;
      RECT 91.02 335.705 91.22 336.435 ;
      RECT 93.21 0.52 93.47 5.16 ;
      RECT 92.69 4.9 93.47 5.16 ;
      RECT 92.69 4.9 92.95 6.64 ;
      RECT 91.84 335.705 92.04 336.435 ;
      RECT 92.335 335.705 92.535 336.435 ;
      RECT 92.835 335.705 93.035 336.435 ;
      RECT 93.335 335.705 93.535 336.435 ;
      RECT 93.83 335.705 94.03 336.435 ;
      RECT 94.575 0.17 95.345 0.94 ;
      RECT 94.575 0.17 94.835 12.9 ;
      RECT 95.085 0.17 95.345 12.9 ;
      RECT 94.065 0.52 94.325 5.815 ;
      RECT 94.65 335.705 94.85 336.435 ;
      RECT 95.595 0.17 96.365 0.43 ;
      RECT 95.595 0.17 95.855 11.5 ;
      RECT 96.105 0.17 96.365 11.5 ;
      RECT 95.145 335.705 95.345 336.435 ;
      RECT 95.645 335.705 95.845 336.435 ;
      RECT 96.145 335.705 96.345 336.435 ;
      RECT 97.635 0.17 98.405 0.43 ;
      RECT 97.635 0.17 97.895 10.48 ;
      RECT 98.145 0.17 98.405 10.99 ;
      RECT 96.64 335.705 96.84 336.435 ;
      RECT 97.46 335.705 97.66 336.435 ;
      RECT 98.655 0.17 99.425 0.94 ;
      RECT 98.655 0.17 98.915 8.7 ;
      RECT 99.165 0.17 99.425 12.9 ;
      RECT 97.955 335.705 98.155 336.435 ;
      RECT 98.455 335.705 98.655 336.435 ;
      RECT 98.955 335.705 99.155 336.435 ;
      RECT 99.45 335.705 99.65 336.435 ;
      RECT 99.675 0.52 99.935 2.485 ;
      RECT 100.27 335.705 100.47 336.435 ;
      RECT 100.54 0.52 100.8 14.11 ;
      RECT 100.765 335.705 100.965 336.435 ;
      RECT 101.05 0.52 101.31 2.335 ;
      RECT 101.265 335.705 101.465 336.435 ;
      RECT 101.765 335.705 101.965 336.435 ;
      RECT 102.26 335.705 102.46 336.435 ;
      RECT 104.45 0.52 104.71 5.16 ;
      RECT 103.93 4.9 104.71 5.16 ;
      RECT 103.93 4.9 104.19 6.64 ;
      RECT 103.08 335.705 103.28 336.435 ;
      RECT 103.575 335.705 103.775 336.435 ;
      RECT 104.075 335.705 104.275 336.435 ;
      RECT 104.575 335.705 104.775 336.435 ;
      RECT 105.07 335.705 105.27 336.435 ;
      RECT 105.815 0.17 106.585 0.94 ;
      RECT 105.815 0.17 106.075 12.9 ;
      RECT 106.325 0.17 106.585 12.9 ;
      RECT 105.305 0.52 105.565 5.815 ;
      RECT 105.89 335.705 106.09 336.435 ;
      RECT 106.835 0.17 107.605 0.43 ;
      RECT 106.835 0.17 107.095 11.5 ;
      RECT 107.345 0.17 107.605 11.5 ;
      RECT 106.385 335.705 106.585 336.435 ;
      RECT 106.885 335.705 107.085 336.435 ;
      RECT 107.385 335.705 107.585 336.435 ;
      RECT 108.875 0.17 109.645 0.43 ;
      RECT 108.875 0.17 109.135 10.48 ;
      RECT 109.385 0.17 109.645 10.99 ;
      RECT 107.88 335.705 108.08 336.435 ;
      RECT 108.7 335.705 108.9 336.435 ;
      RECT 109.895 0.17 110.665 0.94 ;
      RECT 109.895 0.17 110.155 8.7 ;
      RECT 110.405 0.17 110.665 12.9 ;
      RECT 109.195 335.705 109.395 336.435 ;
      RECT 109.695 335.705 109.895 336.435 ;
      RECT 110.195 335.705 110.395 336.435 ;
      RECT 110.69 335.705 110.89 336.435 ;
      RECT 110.915 0.52 111.175 2.485 ;
      RECT 111.51 335.705 111.71 336.435 ;
      RECT 111.78 0.52 112.04 14.11 ;
      RECT 112.005 335.705 112.205 336.435 ;
      RECT 112.29 0.52 112.55 2.335 ;
      RECT 112.505 335.705 112.705 336.435 ;
      RECT 113.005 335.705 113.205 336.435 ;
      RECT 113.5 335.705 113.7 336.435 ;
      RECT 115.69 0.52 115.95 5.16 ;
      RECT 115.17 4.9 115.95 5.16 ;
      RECT 115.17 4.9 115.43 6.64 ;
      RECT 114.32 335.705 114.52 336.435 ;
      RECT 114.815 335.705 115.015 336.435 ;
      RECT 115.315 335.705 115.515 336.435 ;
      RECT 115.815 335.705 116.015 336.435 ;
      RECT 116.31 335.705 116.51 336.435 ;
      RECT 117.055 0.17 117.825 0.94 ;
      RECT 117.055 0.17 117.315 12.9 ;
      RECT 117.565 0.17 117.825 12.9 ;
      RECT 116.545 0.52 116.805 5.815 ;
      RECT 117.13 335.705 117.33 336.435 ;
      RECT 118.075 0.17 118.845 0.43 ;
      RECT 118.075 0.17 118.335 11.5 ;
      RECT 118.585 0.17 118.845 11.5 ;
      RECT 117.625 335.705 117.825 336.435 ;
      RECT 118.125 335.705 118.325 336.435 ;
      RECT 118.625 335.705 118.825 336.435 ;
      RECT 120.115 0.17 120.885 0.43 ;
      RECT 120.115 0.17 120.375 10.48 ;
      RECT 120.625 0.17 120.885 10.99 ;
      RECT 119.12 335.705 119.32 336.435 ;
      RECT 119.94 335.705 120.14 336.435 ;
      RECT 121.135 0.17 121.905 0.94 ;
      RECT 121.135 0.17 121.395 8.7 ;
      RECT 121.645 0.17 121.905 12.9 ;
      RECT 120.435 335.705 120.635 336.435 ;
      RECT 120.935 335.705 121.135 336.435 ;
      RECT 121.435 335.705 121.635 336.435 ;
      RECT 121.93 335.705 122.13 336.435 ;
      RECT 122.155 0.52 122.415 2.485 ;
      RECT 122.75 335.705 122.95 336.435 ;
      RECT 123.02 0.52 123.28 14.11 ;
      RECT 123.245 335.705 123.445 336.435 ;
      RECT 123.53 0.52 123.79 2.335 ;
      RECT 123.745 335.705 123.945 336.435 ;
      RECT 124.245 335.705 124.445 336.435 ;
      RECT 124.74 335.705 124.94 336.435 ;
      RECT 126.93 0.52 127.19 5.16 ;
      RECT 126.41 4.9 127.19 5.16 ;
      RECT 126.41 4.9 126.67 6.64 ;
      RECT 125.56 335.705 125.76 336.435 ;
      RECT 126.055 335.705 126.255 336.435 ;
      RECT 126.555 335.705 126.755 336.435 ;
      RECT 127.055 335.705 127.255 336.435 ;
      RECT 127.55 335.705 127.75 336.435 ;
      RECT 128.295 0.17 129.065 0.94 ;
      RECT 128.295 0.17 128.555 12.9 ;
      RECT 128.805 0.17 129.065 12.9 ;
      RECT 127.785 0.52 128.045 5.815 ;
      RECT 128.37 335.705 128.57 336.435 ;
      RECT 129.315 0.17 130.085 0.43 ;
      RECT 129.315 0.17 129.575 11.5 ;
      RECT 129.825 0.17 130.085 11.5 ;
      RECT 128.865 335.705 129.065 336.435 ;
      RECT 129.365 335.705 129.565 336.435 ;
      RECT 129.865 335.705 130.065 336.435 ;
      RECT 131.355 0.17 132.125 0.43 ;
      RECT 131.355 0.17 131.615 10.48 ;
      RECT 131.865 0.17 132.125 10.99 ;
      RECT 130.36 335.705 130.56 336.435 ;
      RECT 131.18 335.705 131.38 336.435 ;
      RECT 132.375 0.17 133.145 0.94 ;
      RECT 132.375 0.17 132.635 8.7 ;
      RECT 132.885 0.17 133.145 12.9 ;
      RECT 131.675 335.705 131.875 336.435 ;
      RECT 132.175 335.705 132.375 336.435 ;
      RECT 132.675 335.705 132.875 336.435 ;
      RECT 133.17 335.705 133.37 336.435 ;
      RECT 133.395 0.52 133.655 2.485 ;
      RECT 133.99 335.705 134.19 336.435 ;
      RECT 134.26 0.52 134.52 14.11 ;
      RECT 134.485 335.705 134.685 336.435 ;
      RECT 134.77 0.52 135.03 2.335 ;
      RECT 134.985 335.705 135.185 336.435 ;
      RECT 135.485 335.705 135.685 336.435 ;
      RECT 135.98 335.705 136.18 336.435 ;
      RECT 138.17 0.52 138.43 5.16 ;
      RECT 137.65 4.9 138.43 5.16 ;
      RECT 137.65 4.9 137.91 6.64 ;
      RECT 136.8 335.705 137 336.435 ;
      RECT 137.295 335.705 137.495 336.435 ;
      RECT 137.795 335.705 137.995 336.435 ;
      RECT 138.295 335.705 138.495 336.435 ;
      RECT 138.79 335.705 138.99 336.435 ;
      RECT 139.535 0.17 140.305 0.94 ;
      RECT 139.535 0.17 139.795 12.9 ;
      RECT 140.045 0.17 140.305 12.9 ;
      RECT 139.025 0.52 139.285 5.815 ;
      RECT 139.61 335.705 139.81 336.435 ;
      RECT 140.555 0.17 141.325 0.43 ;
      RECT 140.555 0.17 140.815 11.5 ;
      RECT 141.065 0.17 141.325 11.5 ;
      RECT 140.105 335.705 140.305 336.435 ;
      RECT 140.605 335.705 140.805 336.435 ;
      RECT 141.105 335.705 141.305 336.435 ;
      RECT 142.595 0.17 143.365 0.43 ;
      RECT 142.595 0.17 142.855 10.48 ;
      RECT 143.105 0.17 143.365 10.99 ;
      RECT 141.6 335.705 141.8 336.435 ;
      RECT 142.42 335.705 142.62 336.435 ;
      RECT 143.615 0.17 144.385 0.94 ;
      RECT 143.615 0.17 143.875 8.7 ;
      RECT 144.125 0.17 144.385 12.9 ;
      RECT 142.915 335.705 143.115 336.435 ;
      RECT 143.415 335.705 143.615 336.435 ;
      RECT 143.915 335.705 144.115 336.435 ;
      RECT 144.41 335.705 144.61 336.435 ;
      RECT 144.635 0.52 144.895 2.485 ;
      RECT 145.23 335.705 145.43 336.435 ;
      RECT 145.5 0.52 145.76 14.11 ;
      RECT 145.725 335.705 145.925 336.435 ;
      RECT 146.01 0.52 146.27 2.335 ;
      RECT 146.225 335.705 146.425 336.435 ;
      RECT 146.725 335.705 146.925 336.435 ;
      RECT 147.22 335.705 147.42 336.435 ;
      RECT 149.41 0.52 149.67 5.16 ;
      RECT 148.89 4.9 149.67 5.16 ;
      RECT 148.89 4.9 149.15 6.64 ;
      RECT 148.04 335.705 148.24 336.435 ;
      RECT 148.535 335.705 148.735 336.435 ;
      RECT 149.035 335.705 149.235 336.435 ;
      RECT 149.535 335.705 149.735 336.435 ;
      RECT 150.03 335.705 150.23 336.435 ;
      RECT 150.775 0.17 151.545 0.94 ;
      RECT 150.775 0.17 151.035 12.9 ;
      RECT 151.285 0.17 151.545 12.9 ;
      RECT 150.265 0.52 150.525 5.815 ;
      RECT 150.85 335.705 151.05 336.435 ;
      RECT 151.795 0.17 152.565 0.43 ;
      RECT 151.795 0.17 152.055 11.5 ;
      RECT 152.305 0.17 152.565 11.5 ;
      RECT 151.345 335.705 151.545 336.435 ;
      RECT 151.845 335.705 152.045 336.435 ;
      RECT 152.345 335.705 152.545 336.435 ;
      RECT 153.835 0.17 154.605 0.43 ;
      RECT 153.835 0.17 154.095 10.48 ;
      RECT 154.345 0.17 154.605 10.99 ;
      RECT 152.84 335.705 153.04 336.435 ;
      RECT 153.66 335.705 153.86 336.435 ;
      RECT 154.855 0.17 155.625 0.94 ;
      RECT 154.855 0.17 155.115 8.7 ;
      RECT 155.365 0.17 155.625 12.9 ;
      RECT 154.155 335.705 154.355 336.435 ;
      RECT 154.655 335.705 154.855 336.435 ;
      RECT 155.155 335.705 155.355 336.435 ;
      RECT 155.65 335.705 155.85 336.435 ;
      RECT 155.875 0.52 156.135 2.485 ;
      RECT 156.47 335.705 156.67 336.435 ;
      RECT 156.74 0.52 157 14.11 ;
      RECT 156.965 335.705 157.165 336.435 ;
      RECT 157.25 0.52 157.51 2.335 ;
      RECT 157.465 335.705 157.665 336.435 ;
      RECT 157.965 335.705 158.165 336.435 ;
      RECT 158.46 335.705 158.66 336.435 ;
      RECT 160.65 0.52 160.91 5.16 ;
      RECT 160.13 4.9 160.91 5.16 ;
      RECT 160.13 4.9 160.39 6.64 ;
      RECT 159.28 335.705 159.48 336.435 ;
      RECT 159.775 335.705 159.975 336.435 ;
      RECT 160.275 335.705 160.475 336.435 ;
      RECT 160.775 335.705 160.975 336.435 ;
      RECT 161.27 335.705 161.47 336.435 ;
      RECT 162.015 0.17 162.785 0.94 ;
      RECT 162.015 0.17 162.275 12.9 ;
      RECT 162.525 0.17 162.785 12.9 ;
      RECT 161.505 0.52 161.765 5.815 ;
      RECT 162.09 335.705 162.29 336.435 ;
      RECT 163.035 0.17 163.805 0.43 ;
      RECT 163.035 0.17 163.295 11.5 ;
      RECT 163.545 0.17 163.805 11.5 ;
      RECT 162.585 335.705 162.785 336.435 ;
      RECT 163.085 335.705 163.285 336.435 ;
      RECT 163.585 335.705 163.785 336.435 ;
      RECT 165.075 0.17 165.845 0.43 ;
      RECT 165.075 0.17 165.335 10.48 ;
      RECT 165.585 0.17 165.845 10.99 ;
      RECT 164.08 335.705 164.28 336.435 ;
      RECT 164.9 335.705 165.1 336.435 ;
      RECT 166.095 0.17 166.865 0.94 ;
      RECT 166.095 0.17 166.355 8.7 ;
      RECT 166.605 0.17 166.865 12.9 ;
      RECT 165.395 335.705 165.595 336.435 ;
      RECT 165.895 335.705 166.095 336.435 ;
      RECT 166.395 335.705 166.595 336.435 ;
      RECT 166.89 335.705 167.09 336.435 ;
      RECT 167.115 0.52 167.375 2.485 ;
      RECT 167.71 335.705 167.91 336.435 ;
      RECT 167.98 0.52 168.24 14.11 ;
      RECT 168.205 335.705 168.405 336.435 ;
      RECT 168.49 0.52 168.75 2.335 ;
      RECT 168.705 335.705 168.905 336.435 ;
      RECT 169.205 335.705 169.405 336.435 ;
      RECT 169.7 335.705 169.9 336.435 ;
      RECT 171.89 0.52 172.15 5.16 ;
      RECT 171.37 4.9 172.15 5.16 ;
      RECT 171.37 4.9 171.63 6.64 ;
      RECT 170.52 335.705 170.72 336.435 ;
      RECT 171.015 335.705 171.215 336.435 ;
      RECT 171.515 335.705 171.715 336.435 ;
      RECT 172.015 335.705 172.215 336.435 ;
      RECT 172.51 335.705 172.71 336.435 ;
      RECT 173.255 0.17 174.025 0.94 ;
      RECT 173.255 0.17 173.515 12.9 ;
      RECT 173.765 0.17 174.025 12.9 ;
      RECT 172.745 0.52 173.005 5.815 ;
      RECT 173.33 335.705 173.53 336.435 ;
      RECT 174.275 0.17 175.045 0.43 ;
      RECT 174.275 0.17 174.535 11.5 ;
      RECT 174.785 0.17 175.045 11.5 ;
      RECT 173.825 335.705 174.025 336.435 ;
      RECT 174.325 335.705 174.525 336.435 ;
      RECT 174.825 335.705 175.025 336.435 ;
      RECT 176.315 0.17 177.085 0.43 ;
      RECT 176.315 0.17 176.575 10.48 ;
      RECT 176.825 0.17 177.085 10.99 ;
      RECT 175.32 335.705 175.52 336.435 ;
      RECT 176.14 335.705 176.34 336.435 ;
      RECT 177.335 0.17 178.105 0.94 ;
      RECT 177.335 0.17 177.595 8.7 ;
      RECT 177.845 0.17 178.105 12.9 ;
      RECT 176.635 335.705 176.835 336.435 ;
      RECT 177.135 335.705 177.335 336.435 ;
      RECT 177.635 335.705 177.835 336.435 ;
      RECT 178.13 335.705 178.33 336.435 ;
      RECT 178.355 0.52 178.615 2.485 ;
      RECT 178.95 335.705 179.15 336.435 ;
      RECT 179.22 0.52 179.48 14.11 ;
      RECT 179.445 335.705 179.645 336.435 ;
      RECT 179.73 0.52 179.99 2.335 ;
      RECT 179.945 335.705 180.145 336.435 ;
      RECT 180.445 335.705 180.645 336.435 ;
      RECT 182.435 0.17 183.205 0.43 ;
      RECT 182.435 0.17 182.695 8.7 ;
      RECT 182.945 0.17 183.205 8.7 ;
      RECT 183.455 0.17 184.225 0.94 ;
      RECT 183.455 0.17 183.715 8.7 ;
      RECT 183.965 0.17 184.225 8.7 ;
      RECT 184.475 0.17 185.245 0.43 ;
      RECT 184.475 0.17 184.735 8.7 ;
      RECT 184.985 0.17 185.245 8.7 ;
      RECT 185.495 0.17 186.265 0.94 ;
      RECT 185.495 0.17 185.755 8.7 ;
      RECT 186.005 0.17 186.265 8.7 ;
      RECT 186.515 0.17 187.285 0.43 ;
      RECT 186.515 0.17 186.775 8.7 ;
      RECT 187.025 0.17 187.285 8.7 ;
      RECT 187.535 0.17 188.305 0.94 ;
      RECT 187.535 0.17 187.795 8.7 ;
      RECT 188.045 0.17 188.305 8.7 ;
      RECT 180.94 335.705 181.14 336.435 ;
      RECT 181.76 335.705 181.96 336.435 ;
      RECT 182.755 335.705 182.955 336.435 ;
      RECT 190.24 0.17 191.01 0.94 ;
      RECT 190.24 0.17 190.5 8.7 ;
      RECT 190.75 0.17 191.01 8.7 ;
      RECT 188.71 0.3 188.97 8.7 ;
      RECT 189.22 0 189.48 8.7 ;
      RECT 189.73 0 189.99 8.7 ;
      RECT 191.26 0 191.52 8.7 ;
      RECT 191.77 0 192.03 8.7 ;
      RECT 192.28 0.52 192.54 8.7 ;
      RECT 192.79 0.52 193.05 8.7 ;
      RECT 193.3 0.52 193.56 8.7 ;
      RECT 195.34 0.17 196.11 0.94 ;
      RECT 195.34 0.17 195.6 8.7 ;
      RECT 195.85 0.17 196.11 8.7 ;
      RECT 196.36 0.17 197.13 0.43 ;
      RECT 196.36 0.17 196.62 8.7 ;
      RECT 196.87 0.17 197.13 8.7 ;
      RECT 193.81 0.52 194.07 8.7 ;
      RECT 194.32 0 194.58 8.7 ;
      RECT 194.83 0 195.09 8.7 ;
      RECT 197.38 0.3 197.64 8.7 ;
      RECT 197.89 0.3 198.15 8.7 ;
      RECT 199.93 0.17 200.7 0.94 ;
      RECT 199.93 0.17 200.19 8.7 ;
      RECT 200.44 0.17 200.7 8.7 ;
      RECT 198.4 0.3 198.66 8.7 ;
      RECT 198.91 0.3 199.17 8.7 ;
      RECT 199.42 0.3 199.68 8.7 ;
      RECT 200.95 0.52 201.21 8.7 ;
      RECT 201.46 0.52 201.72 8.7 ;
      RECT 201.97 0.3 202.23 8.7 ;
      RECT 202.48 0.52 202.74 8.7 ;
      RECT 202.99 0.52 203.25 8.7 ;
      RECT 203.5 0.3 203.76 8.7 ;
      RECT 204.01 0.52 204.27 8.7 ;
      RECT 204.52 0.52 204.78 8.7 ;
      RECT 205.03 0.52 205.29 8.7 ;
      RECT 205.54 0.52 205.8 8.7 ;
      RECT 206.05 0.52 206.31 8.7 ;
      RECT 206.56 0.3 206.82 8.7 ;
      RECT 207.07 0.52 207.33 8.7 ;
      RECT 207.58 0.52 207.84 8.7 ;
      RECT 208.09 0.3 208.35 8.7 ;
      RECT 210.13 0.17 210.9 0.94 ;
      RECT 210.13 0.17 210.39 8.7 ;
      RECT 210.64 0.17 210.9 8.7 ;
      RECT 208.6 0.52 208.86 8.7 ;
      RECT 209.11 0.52 209.37 8.7 ;
      RECT 209.62 0.3 209.88 8.7 ;
      RECT 211.15 0.52 211.41 8.7 ;
      RECT 211.66 0.52 211.92 8.7 ;
      RECT 212.17 0.52 212.43 8.7 ;
      RECT 212.68 0.52 212.94 8.7 ;
      RECT 213.19 0.52 213.45 8.7 ;
      RECT 213.7 0.52 213.96 8.7 ;
      RECT 214.21 0.52 214.47 8.7 ;
      RECT 216.25 0.17 217.02 0.94 ;
      RECT 216.25 0.17 216.51 8.7 ;
      RECT 216.76 0.17 217.02 8.7 ;
      RECT 214.72 0.52 214.98 8.7 ;
      RECT 215.23 0 215.49 8.7 ;
      RECT 215.74 0 216 8.7 ;
      RECT 217.27 0.52 217.53 8.7 ;
      RECT 219.31 0.17 220.08 0.43 ;
      RECT 219.31 0.17 219.57 8.7 ;
      RECT 219.82 0.17 220.08 8.7 ;
      RECT 217.78 0.52 218.04 8.7 ;
      RECT 218.29 0.3 218.55 8.7 ;
      RECT 218.8 0.3 219.06 8.7 ;
      RECT 220.33 0.3 220.59 8.7 ;
      RECT 220.84 0.3 221.1 8.7 ;
      RECT 221.35 0.3 221.61 8.7 ;
      RECT 221.86 0.3 222.12 8.7 ;
      RECT 222.37 0.52 222.63 8.7 ;
      RECT 222.88 0.52 223.14 8.7 ;
      RECT 224.92 0.17 225.69 0.43 ;
      RECT 224.92 0.17 225.18 8.7 ;
      RECT 225.43 0.17 225.69 8.7 ;
      RECT 225.94 0.17 226.71 0.94 ;
      RECT 225.94 0.17 226.2 25.5 ;
      RECT 226.45 0.17 226.71 33.9 ;
      RECT 226.96 0.17 227.73 0.43 ;
      RECT 226.96 0.17 227.22 8.7 ;
      RECT 227.47 0.17 227.73 8.7 ;
      RECT 228.335 0.17 229.105 0.94 ;
      RECT 228.335 0.17 228.595 8.7 ;
      RECT 228.845 0.17 229.105 8.7 ;
      RECT 229.355 0.17 230.125 0.43 ;
      RECT 229.355 0.17 229.615 8.7 ;
      RECT 229.865 0.17 230.125 8.7 ;
      RECT 230.375 0.17 231.145 0.94 ;
      RECT 230.375 0.17 230.635 8.7 ;
      RECT 230.885 0.17 231.145 8.7 ;
      RECT 231.395 0.17 232.165 0.43 ;
      RECT 231.395 0.17 231.655 8.7 ;
      RECT 231.905 0.17 232.165 8.7 ;
      RECT 232.415 0.17 233.185 0.94 ;
      RECT 232.415 0.17 232.675 8.7 ;
      RECT 232.925 0.17 233.185 8.7 ;
      RECT 223.39 0.3 223.65 8.7 ;
      RECT 233.435 0.17 234.205 0.43 ;
      RECT 233.435 0.17 233.695 8.7 ;
      RECT 233.945 0.17 234.205 8.7 ;
      RECT 223.9 0.3 224.16 8.7 ;
      RECT 224.41 0.52 224.67 8.7 ;
      RECT 233.685 335.705 233.885 336.435 ;
      RECT 234.68 335.705 234.88 336.435 ;
      RECT 235.5 335.705 235.7 336.435 ;
      RECT 235.995 335.705 236.195 336.435 ;
      RECT 236.495 335.705 236.695 336.435 ;
      RECT 236.65 0.52 236.91 2.335 ;
      RECT 236.995 335.705 237.195 336.435 ;
      RECT 237.16 0.52 237.42 14.11 ;
      RECT 237.49 335.705 237.69 336.435 ;
      RECT 238.535 0.17 239.305 0.94 ;
      RECT 239.045 0.17 239.305 8.7 ;
      RECT 238.535 0.17 238.795 12.9 ;
      RECT 238.025 0.52 238.285 2.485 ;
      RECT 238.31 335.705 238.51 336.435 ;
      RECT 239.555 0.17 240.325 0.43 ;
      RECT 240.065 0.17 240.325 10.48 ;
      RECT 239.555 0.17 239.815 10.99 ;
      RECT 238.805 335.705 239.005 336.435 ;
      RECT 239.305 335.705 239.505 336.435 ;
      RECT 239.805 335.705 240.005 336.435 ;
      RECT 240.3 335.705 240.5 336.435 ;
      RECT 241.595 0.17 242.365 0.43 ;
      RECT 241.595 0.17 241.855 11.5 ;
      RECT 242.105 0.17 242.365 11.5 ;
      RECT 241.12 335.705 241.32 336.435 ;
      RECT 241.615 335.705 241.815 336.435 ;
      RECT 242.615 0.17 243.385 0.94 ;
      RECT 242.615 0.17 242.875 12.9 ;
      RECT 243.125 0.17 243.385 12.9 ;
      RECT 242.115 335.705 242.315 336.435 ;
      RECT 242.615 335.705 242.815 336.435 ;
      RECT 243.11 335.705 243.31 336.435 ;
      RECT 243.635 0.52 243.895 5.815 ;
      RECT 244.49 0.52 244.75 5.16 ;
      RECT 244.49 4.9 245.27 5.16 ;
      RECT 245.01 4.9 245.27 6.64 ;
      RECT 243.93 335.705 244.13 336.435 ;
      RECT 244.425 335.705 244.625 336.435 ;
      RECT 244.925 335.705 245.125 336.435 ;
      RECT 245.425 335.705 245.625 336.435 ;
      RECT 245.92 335.705 246.12 336.435 ;
      RECT 246.74 335.705 246.94 336.435 ;
      RECT 247.235 335.705 247.435 336.435 ;
      RECT 247.735 335.705 247.935 336.435 ;
      RECT 247.89 0.52 248.15 2.335 ;
      RECT 248.235 335.705 248.435 336.435 ;
      RECT 248.4 0.52 248.66 14.11 ;
      RECT 248.73 335.705 248.93 336.435 ;
      RECT 249.775 0.17 250.545 0.94 ;
      RECT 250.285 0.17 250.545 8.7 ;
      RECT 249.775 0.17 250.035 12.9 ;
      RECT 249.265 0.52 249.525 2.485 ;
      RECT 249.55 335.705 249.75 336.435 ;
      RECT 250.795 0.17 251.565 0.43 ;
      RECT 251.305 0.17 251.565 10.48 ;
      RECT 250.795 0.17 251.055 10.99 ;
      RECT 250.045 335.705 250.245 336.435 ;
      RECT 250.545 335.705 250.745 336.435 ;
      RECT 251.045 335.705 251.245 336.435 ;
      RECT 251.54 335.705 251.74 336.435 ;
      RECT 252.835 0.17 253.605 0.43 ;
      RECT 252.835 0.17 253.095 11.5 ;
      RECT 253.345 0.17 253.605 11.5 ;
      RECT 252.36 335.705 252.56 336.435 ;
      RECT 252.855 335.705 253.055 336.435 ;
      RECT 253.855 0.17 254.625 0.94 ;
      RECT 253.855 0.17 254.115 12.9 ;
      RECT 254.365 0.17 254.625 12.9 ;
      RECT 253.355 335.705 253.555 336.435 ;
      RECT 253.855 335.705 254.055 336.435 ;
      RECT 254.35 335.705 254.55 336.435 ;
      RECT 254.875 0.52 255.135 5.815 ;
      RECT 255.73 0.52 255.99 5.16 ;
      RECT 255.73 4.9 256.51 5.16 ;
      RECT 256.25 4.9 256.51 6.64 ;
      RECT 255.17 335.705 255.37 336.435 ;
      RECT 255.665 335.705 255.865 336.435 ;
      RECT 256.165 335.705 256.365 336.435 ;
      RECT 256.665 335.705 256.865 336.435 ;
      RECT 257.16 335.705 257.36 336.435 ;
      RECT 257.98 335.705 258.18 336.435 ;
      RECT 258.475 335.705 258.675 336.435 ;
      RECT 258.975 335.705 259.175 336.435 ;
      RECT 259.13 0.52 259.39 2.335 ;
      RECT 259.475 335.705 259.675 336.435 ;
      RECT 259.64 0.52 259.9 14.11 ;
      RECT 259.97 335.705 260.17 336.435 ;
      RECT 261.015 0.17 261.785 0.94 ;
      RECT 261.525 0.17 261.785 8.7 ;
      RECT 261.015 0.17 261.275 12.9 ;
      RECT 260.505 0.52 260.765 2.485 ;
      RECT 260.79 335.705 260.99 336.435 ;
      RECT 262.035 0.17 262.805 0.43 ;
      RECT 262.545 0.17 262.805 10.48 ;
      RECT 262.035 0.17 262.295 10.99 ;
      RECT 261.285 335.705 261.485 336.435 ;
      RECT 261.785 335.705 261.985 336.435 ;
      RECT 262.285 335.705 262.485 336.435 ;
      RECT 262.78 335.705 262.98 336.435 ;
      RECT 264.075 0.17 264.845 0.43 ;
      RECT 264.075 0.17 264.335 11.5 ;
      RECT 264.585 0.17 264.845 11.5 ;
      RECT 263.6 335.705 263.8 336.435 ;
      RECT 264.095 335.705 264.295 336.435 ;
      RECT 265.095 0.17 265.865 0.94 ;
      RECT 265.095 0.17 265.355 12.9 ;
      RECT 265.605 0.17 265.865 12.9 ;
      RECT 264.595 335.705 264.795 336.435 ;
      RECT 265.095 335.705 265.295 336.435 ;
      RECT 265.59 335.705 265.79 336.435 ;
      RECT 266.115 0.52 266.375 5.815 ;
      RECT 266.97 0.52 267.23 5.16 ;
      RECT 266.97 4.9 267.75 5.16 ;
      RECT 267.49 4.9 267.75 6.64 ;
      RECT 266.41 335.705 266.61 336.435 ;
      RECT 266.905 335.705 267.105 336.435 ;
      RECT 267.405 335.705 267.605 336.435 ;
      RECT 267.905 335.705 268.105 336.435 ;
      RECT 268.4 335.705 268.6 336.435 ;
      RECT 269.22 335.705 269.42 336.435 ;
      RECT 269.715 335.705 269.915 336.435 ;
      RECT 270.215 335.705 270.415 336.435 ;
      RECT 270.37 0.52 270.63 2.335 ;
      RECT 270.715 335.705 270.915 336.435 ;
      RECT 270.88 0.52 271.14 14.11 ;
      RECT 271.21 335.705 271.41 336.435 ;
      RECT 272.255 0.17 273.025 0.94 ;
      RECT 272.765 0.17 273.025 8.7 ;
      RECT 272.255 0.17 272.515 12.9 ;
      RECT 271.745 0.52 272.005 2.485 ;
      RECT 272.03 335.705 272.23 336.435 ;
      RECT 273.275 0.17 274.045 0.43 ;
      RECT 273.785 0.17 274.045 10.48 ;
      RECT 273.275 0.17 273.535 10.99 ;
      RECT 272.525 335.705 272.725 336.435 ;
      RECT 273.025 335.705 273.225 336.435 ;
      RECT 273.525 335.705 273.725 336.435 ;
      RECT 274.02 335.705 274.22 336.435 ;
      RECT 275.315 0.17 276.085 0.43 ;
      RECT 275.315 0.17 275.575 11.5 ;
      RECT 275.825 0.17 276.085 11.5 ;
      RECT 274.84 335.705 275.04 336.435 ;
      RECT 275.335 335.705 275.535 336.435 ;
      RECT 276.335 0.17 277.105 0.94 ;
      RECT 276.335 0.17 276.595 12.9 ;
      RECT 276.845 0.17 277.105 12.9 ;
      RECT 275.835 335.705 276.035 336.435 ;
      RECT 276.335 335.705 276.535 336.435 ;
      RECT 276.83 335.705 277.03 336.435 ;
      RECT 277.355 0.52 277.615 5.815 ;
      RECT 278.21 0.52 278.47 5.16 ;
      RECT 278.21 4.9 278.99 5.16 ;
      RECT 278.73 4.9 278.99 6.64 ;
      RECT 277.65 335.705 277.85 336.435 ;
      RECT 278.145 335.705 278.345 336.435 ;
      RECT 278.645 335.705 278.845 336.435 ;
      RECT 279.145 335.705 279.345 336.435 ;
      RECT 279.64 335.705 279.84 336.435 ;
      RECT 280.46 335.705 280.66 336.435 ;
      RECT 280.955 335.705 281.155 336.435 ;
      RECT 281.455 335.705 281.655 336.435 ;
      RECT 281.61 0.52 281.87 2.335 ;
      RECT 281.955 335.705 282.155 336.435 ;
      RECT 282.12 0.52 282.38 14.11 ;
      RECT 282.45 335.705 282.65 336.435 ;
      RECT 283.495 0.17 284.265 0.94 ;
      RECT 284.005 0.17 284.265 8.7 ;
      RECT 283.495 0.17 283.755 12.9 ;
      RECT 282.985 0.52 283.245 2.485 ;
      RECT 283.27 335.705 283.47 336.435 ;
      RECT 284.515 0.17 285.285 0.43 ;
      RECT 285.025 0.17 285.285 10.48 ;
      RECT 284.515 0.17 284.775 10.99 ;
      RECT 283.765 335.705 283.965 336.435 ;
      RECT 284.265 335.705 284.465 336.435 ;
      RECT 284.765 335.705 284.965 336.435 ;
      RECT 285.26 335.705 285.46 336.435 ;
      RECT 286.555 0.17 287.325 0.43 ;
      RECT 286.555 0.17 286.815 11.5 ;
      RECT 287.065 0.17 287.325 11.5 ;
      RECT 286.08 335.705 286.28 336.435 ;
      RECT 286.575 335.705 286.775 336.435 ;
      RECT 287.575 0.17 288.345 0.94 ;
      RECT 287.575 0.17 287.835 12.9 ;
      RECT 288.085 0.17 288.345 12.9 ;
      RECT 287.075 335.705 287.275 336.435 ;
      RECT 287.575 335.705 287.775 336.435 ;
      RECT 288.07 335.705 288.27 336.435 ;
      RECT 288.595 0.52 288.855 5.815 ;
      RECT 289.45 0.52 289.71 5.16 ;
      RECT 289.45 4.9 290.23 5.16 ;
      RECT 289.97 4.9 290.23 6.64 ;
      RECT 288.89 335.705 289.09 336.435 ;
      RECT 289.385 335.705 289.585 336.435 ;
      RECT 289.885 335.705 290.085 336.435 ;
      RECT 290.385 335.705 290.585 336.435 ;
      RECT 290.88 335.705 291.08 336.435 ;
      RECT 291.7 335.705 291.9 336.435 ;
      RECT 292.195 335.705 292.395 336.435 ;
      RECT 292.695 335.705 292.895 336.435 ;
      RECT 292.85 0.52 293.11 2.335 ;
      RECT 293.195 335.705 293.395 336.435 ;
      RECT 293.36 0.52 293.62 14.11 ;
      RECT 293.69 335.705 293.89 336.435 ;
      RECT 294.735 0.17 295.505 0.94 ;
      RECT 295.245 0.17 295.505 8.7 ;
      RECT 294.735 0.17 294.995 12.9 ;
      RECT 294.225 0.52 294.485 2.485 ;
      RECT 294.51 335.705 294.71 336.435 ;
      RECT 295.755 0.17 296.525 0.43 ;
      RECT 296.265 0.17 296.525 10.48 ;
      RECT 295.755 0.17 296.015 10.99 ;
      RECT 295.005 335.705 295.205 336.435 ;
      RECT 295.505 335.705 295.705 336.435 ;
      RECT 296.005 335.705 296.205 336.435 ;
      RECT 296.5 335.705 296.7 336.435 ;
      RECT 297.795 0.17 298.565 0.43 ;
      RECT 297.795 0.17 298.055 11.5 ;
      RECT 298.305 0.17 298.565 11.5 ;
      RECT 297.32 335.705 297.52 336.435 ;
      RECT 297.815 335.705 298.015 336.435 ;
      RECT 298.815 0.17 299.585 0.94 ;
      RECT 298.815 0.17 299.075 12.9 ;
      RECT 299.325 0.17 299.585 12.9 ;
      RECT 298.315 335.705 298.515 336.435 ;
      RECT 298.815 335.705 299.015 336.435 ;
      RECT 299.31 335.705 299.51 336.435 ;
      RECT 299.835 0.52 300.095 5.815 ;
      RECT 300.69 0.52 300.95 5.16 ;
      RECT 300.69 4.9 301.47 5.16 ;
      RECT 301.21 4.9 301.47 6.64 ;
      RECT 300.13 335.705 300.33 336.435 ;
      RECT 300.625 335.705 300.825 336.435 ;
      RECT 301.125 335.705 301.325 336.435 ;
      RECT 301.625 335.705 301.825 336.435 ;
      RECT 302.12 335.705 302.32 336.435 ;
      RECT 302.94 335.705 303.14 336.435 ;
      RECT 303.435 335.705 303.635 336.435 ;
      RECT 303.935 335.705 304.135 336.435 ;
      RECT 304.09 0.52 304.35 2.335 ;
      RECT 304.435 335.705 304.635 336.435 ;
      RECT 304.6 0.52 304.86 14.11 ;
      RECT 304.93 335.705 305.13 336.435 ;
      RECT 305.975 0.17 306.745 0.94 ;
      RECT 306.485 0.17 306.745 8.7 ;
      RECT 305.975 0.17 306.235 12.9 ;
      RECT 305.465 0.52 305.725 2.485 ;
      RECT 305.75 335.705 305.95 336.435 ;
      RECT 306.995 0.17 307.765 0.43 ;
      RECT 307.505 0.17 307.765 10.48 ;
      RECT 306.995 0.17 307.255 10.99 ;
      RECT 306.245 335.705 306.445 336.435 ;
      RECT 306.745 335.705 306.945 336.435 ;
      RECT 307.245 335.705 307.445 336.435 ;
      RECT 307.74 335.705 307.94 336.435 ;
      RECT 309.035 0.17 309.805 0.43 ;
      RECT 309.035 0.17 309.295 11.5 ;
      RECT 309.545 0.17 309.805 11.5 ;
      RECT 308.56 335.705 308.76 336.435 ;
      RECT 309.055 335.705 309.255 336.435 ;
      RECT 310.055 0.17 310.825 0.94 ;
      RECT 310.055 0.17 310.315 12.9 ;
      RECT 310.565 0.17 310.825 12.9 ;
      RECT 309.555 335.705 309.755 336.435 ;
      RECT 310.055 335.705 310.255 336.435 ;
      RECT 310.55 335.705 310.75 336.435 ;
      RECT 311.075 0.52 311.335 5.815 ;
      RECT 311.93 0.52 312.19 5.16 ;
      RECT 311.93 4.9 312.71 5.16 ;
      RECT 312.45 4.9 312.71 6.64 ;
      RECT 311.37 335.705 311.57 336.435 ;
      RECT 311.865 335.705 312.065 336.435 ;
      RECT 312.365 335.705 312.565 336.435 ;
      RECT 312.865 335.705 313.065 336.435 ;
      RECT 313.36 335.705 313.56 336.435 ;
      RECT 314.18 335.705 314.38 336.435 ;
      RECT 314.675 335.705 314.875 336.435 ;
      RECT 315.175 335.705 315.375 336.435 ;
      RECT 315.33 0.52 315.59 2.335 ;
      RECT 315.675 335.705 315.875 336.435 ;
      RECT 315.84 0.52 316.1 14.11 ;
      RECT 316.17 335.705 316.37 336.435 ;
      RECT 317.215 0.17 317.985 0.94 ;
      RECT 317.725 0.17 317.985 8.7 ;
      RECT 317.215 0.17 317.475 12.9 ;
      RECT 316.705 0.52 316.965 2.485 ;
      RECT 316.99 335.705 317.19 336.435 ;
      RECT 318.235 0.17 319.005 0.43 ;
      RECT 318.745 0.17 319.005 10.48 ;
      RECT 318.235 0.17 318.495 10.99 ;
      RECT 317.485 335.705 317.685 336.435 ;
      RECT 317.985 335.705 318.185 336.435 ;
      RECT 318.485 335.705 318.685 336.435 ;
      RECT 318.98 335.705 319.18 336.435 ;
      RECT 320.275 0.17 321.045 0.43 ;
      RECT 320.275 0.17 320.535 11.5 ;
      RECT 320.785 0.17 321.045 11.5 ;
      RECT 319.8 335.705 320 336.435 ;
      RECT 320.295 335.705 320.495 336.435 ;
      RECT 321.295 0.17 322.065 0.94 ;
      RECT 321.295 0.17 321.555 12.9 ;
      RECT 321.805 0.17 322.065 12.9 ;
      RECT 320.795 335.705 320.995 336.435 ;
      RECT 321.295 335.705 321.495 336.435 ;
      RECT 321.79 335.705 321.99 336.435 ;
      RECT 322.315 0.52 322.575 5.815 ;
      RECT 323.17 0.52 323.43 5.16 ;
      RECT 323.17 4.9 323.95 5.16 ;
      RECT 323.69 4.9 323.95 6.64 ;
      RECT 322.61 335.705 322.81 336.435 ;
      RECT 323.105 335.705 323.305 336.435 ;
      RECT 323.605 335.705 323.805 336.435 ;
      RECT 324.105 335.705 324.305 336.435 ;
      RECT 324.6 335.705 324.8 336.435 ;
      RECT 325.42 335.705 325.62 336.435 ;
      RECT 325.915 335.705 326.115 336.435 ;
      RECT 326.415 335.705 326.615 336.435 ;
      RECT 326.57 0.52 326.83 2.335 ;
      RECT 326.915 335.705 327.115 336.435 ;
      RECT 327.08 0.52 327.34 14.11 ;
      RECT 327.41 335.705 327.61 336.435 ;
      RECT 328.455 0.17 329.225 0.94 ;
      RECT 328.965 0.17 329.225 8.7 ;
      RECT 328.455 0.17 328.715 12.9 ;
      RECT 327.945 0.52 328.205 2.485 ;
      RECT 328.23 335.705 328.43 336.435 ;
      RECT 329.475 0.17 330.245 0.43 ;
      RECT 329.985 0.17 330.245 10.48 ;
      RECT 329.475 0.17 329.735 10.99 ;
      RECT 328.725 335.705 328.925 336.435 ;
      RECT 329.225 335.705 329.425 336.435 ;
      RECT 329.725 335.705 329.925 336.435 ;
      RECT 330.22 335.705 330.42 336.435 ;
      RECT 331.515 0.17 332.285 0.43 ;
      RECT 331.515 0.17 331.775 11.5 ;
      RECT 332.025 0.17 332.285 11.5 ;
      RECT 331.04 335.705 331.24 336.435 ;
      RECT 331.535 335.705 331.735 336.435 ;
      RECT 332.535 0.17 333.305 0.94 ;
      RECT 332.535 0.17 332.795 12.9 ;
      RECT 333.045 0.17 333.305 12.9 ;
      RECT 332.035 335.705 332.235 336.435 ;
      RECT 332.535 335.705 332.735 336.435 ;
      RECT 333.03 335.705 333.23 336.435 ;
      RECT 333.555 0.52 333.815 5.815 ;
      RECT 334.41 0.52 334.67 5.16 ;
      RECT 334.41 4.9 335.19 5.16 ;
      RECT 334.93 4.9 335.19 6.64 ;
      RECT 333.85 335.705 334.05 336.435 ;
      RECT 334.345 335.705 334.545 336.435 ;
      RECT 334.845 335.705 335.045 336.435 ;
      RECT 335.345 335.705 335.545 336.435 ;
      RECT 335.84 335.705 336.04 336.435 ;
      RECT 336.66 335.705 336.86 336.435 ;
      RECT 337.155 335.705 337.355 336.435 ;
      RECT 337.655 335.705 337.855 336.435 ;
      RECT 337.81 0.52 338.07 2.335 ;
      RECT 338.155 335.705 338.355 336.435 ;
      RECT 338.32 0.52 338.58 14.11 ;
      RECT 338.65 335.705 338.85 336.435 ;
      RECT 339.695 0.17 340.465 0.94 ;
      RECT 340.205 0.17 340.465 8.7 ;
      RECT 339.695 0.17 339.955 12.9 ;
      RECT 339.185 0.52 339.445 2.485 ;
      RECT 339.47 335.705 339.67 336.435 ;
      RECT 340.715 0.17 341.485 0.43 ;
      RECT 341.225 0.17 341.485 10.48 ;
      RECT 340.715 0.17 340.975 10.99 ;
      RECT 339.965 335.705 340.165 336.435 ;
      RECT 340.465 335.705 340.665 336.435 ;
      RECT 340.965 335.705 341.165 336.435 ;
      RECT 341.46 335.705 341.66 336.435 ;
      RECT 342.755 0.17 343.525 0.43 ;
      RECT 342.755 0.17 343.015 11.5 ;
      RECT 343.265 0.17 343.525 11.5 ;
      RECT 342.28 335.705 342.48 336.435 ;
      RECT 342.775 335.705 342.975 336.435 ;
      RECT 343.775 0.17 344.545 0.94 ;
      RECT 343.775 0.17 344.035 12.9 ;
      RECT 344.285 0.17 344.545 12.9 ;
      RECT 343.275 335.705 343.475 336.435 ;
      RECT 343.775 335.705 343.975 336.435 ;
      RECT 344.27 335.705 344.47 336.435 ;
      RECT 344.795 0.52 345.055 5.815 ;
      RECT 345.65 0.52 345.91 5.16 ;
      RECT 345.65 4.9 346.43 5.16 ;
      RECT 346.17 4.9 346.43 6.64 ;
      RECT 345.09 335.705 345.29 336.435 ;
      RECT 345.585 335.705 345.785 336.435 ;
      RECT 346.085 335.705 346.285 336.435 ;
      RECT 346.585 335.705 346.785 336.435 ;
      RECT 347.08 335.705 347.28 336.435 ;
      RECT 347.9 335.705 348.1 336.435 ;
      RECT 348.395 335.705 348.595 336.435 ;
      RECT 348.895 335.705 349.095 336.435 ;
      RECT 349.05 0.52 349.31 2.335 ;
      RECT 349.395 335.705 349.595 336.435 ;
      RECT 349.56 0.52 349.82 14.11 ;
      RECT 349.89 335.705 350.09 336.435 ;
      RECT 350.935 0.17 351.705 0.94 ;
      RECT 351.445 0.17 351.705 8.7 ;
      RECT 350.935 0.17 351.195 12.9 ;
      RECT 350.425 0.52 350.685 2.485 ;
      RECT 350.71 335.705 350.91 336.435 ;
      RECT 351.955 0.17 352.725 0.43 ;
      RECT 352.465 0.17 352.725 10.48 ;
      RECT 351.955 0.17 352.215 10.99 ;
      RECT 351.205 335.705 351.405 336.435 ;
      RECT 351.705 335.705 351.905 336.435 ;
      RECT 352.205 335.705 352.405 336.435 ;
      RECT 352.7 335.705 352.9 336.435 ;
      RECT 353.995 0.17 354.765 0.43 ;
      RECT 353.995 0.17 354.255 11.5 ;
      RECT 354.505 0.17 354.765 11.5 ;
      RECT 353.52 335.705 353.72 336.435 ;
      RECT 354.015 335.705 354.215 336.435 ;
      RECT 355.015 0.17 355.785 0.94 ;
      RECT 355.015 0.17 355.275 12.9 ;
      RECT 355.525 0.17 355.785 12.9 ;
      RECT 354.515 335.705 354.715 336.435 ;
      RECT 355.015 335.705 355.215 336.435 ;
      RECT 355.51 335.705 355.71 336.435 ;
      RECT 356.035 0.52 356.295 5.815 ;
      RECT 356.89 0.52 357.15 5.16 ;
      RECT 356.89 4.9 357.67 5.16 ;
      RECT 357.41 4.9 357.67 6.64 ;
      RECT 356.33 335.705 356.53 336.435 ;
      RECT 356.825 335.705 357.025 336.435 ;
      RECT 357.325 335.705 357.525 336.435 ;
      RECT 357.825 335.705 358.025 336.435 ;
      RECT 358.32 335.705 358.52 336.435 ;
      RECT 359.14 335.705 359.34 336.435 ;
      RECT 359.635 335.705 359.835 336.435 ;
      RECT 360.135 335.705 360.335 336.435 ;
      RECT 360.29 0.52 360.55 2.335 ;
      RECT 360.635 335.705 360.835 336.435 ;
      RECT 360.8 0.52 361.06 14.11 ;
      RECT 361.13 335.705 361.33 336.435 ;
      RECT 362.175 0.17 362.945 0.94 ;
      RECT 362.685 0.17 362.945 8.7 ;
      RECT 362.175 0.17 362.435 12.9 ;
      RECT 361.665 0.52 361.925 2.485 ;
      RECT 361.95 335.705 362.15 336.435 ;
      RECT 363.195 0.17 363.965 0.43 ;
      RECT 363.705 0.17 363.965 10.48 ;
      RECT 363.195 0.17 363.455 10.99 ;
      RECT 362.445 335.705 362.645 336.435 ;
      RECT 362.945 335.705 363.145 336.435 ;
      RECT 363.445 335.705 363.645 336.435 ;
      RECT 363.94 335.705 364.14 336.435 ;
      RECT 365.235 0.17 366.005 0.43 ;
      RECT 365.235 0.17 365.495 11.5 ;
      RECT 365.745 0.17 366.005 11.5 ;
      RECT 364.76 335.705 364.96 336.435 ;
      RECT 365.255 335.705 365.455 336.435 ;
      RECT 366.255 0.17 367.025 0.94 ;
      RECT 366.255 0.17 366.515 12.9 ;
      RECT 366.765 0.17 367.025 12.9 ;
      RECT 365.755 335.705 365.955 336.435 ;
      RECT 366.255 335.705 366.455 336.435 ;
      RECT 366.75 335.705 366.95 336.435 ;
      RECT 367.275 0.52 367.535 5.815 ;
      RECT 368.13 0.52 368.39 5.16 ;
      RECT 368.13 4.9 368.91 5.16 ;
      RECT 368.65 4.9 368.91 6.64 ;
      RECT 367.57 335.705 367.77 336.435 ;
      RECT 368.065 335.705 368.265 336.435 ;
      RECT 368.565 335.705 368.765 336.435 ;
      RECT 369.065 335.705 369.265 336.435 ;
      RECT 369.56 335.705 369.76 336.435 ;
      RECT 370.38 335.705 370.58 336.435 ;
      RECT 370.875 335.705 371.075 336.435 ;
      RECT 371.375 335.705 371.575 336.435 ;
      RECT 371.53 0.52 371.79 2.335 ;
      RECT 371.875 335.705 372.075 336.435 ;
      RECT 372.04 0.52 372.3 14.11 ;
      RECT 372.37 335.705 372.57 336.435 ;
      RECT 373.415 0.17 374.185 0.94 ;
      RECT 373.925 0.17 374.185 8.7 ;
      RECT 373.415 0.17 373.675 12.9 ;
      RECT 372.905 0.52 373.165 2.485 ;
      RECT 373.19 335.705 373.39 336.435 ;
      RECT 374.435 0.17 375.205 0.43 ;
      RECT 374.945 0.17 375.205 10.48 ;
      RECT 374.435 0.17 374.695 10.99 ;
      RECT 373.685 335.705 373.885 336.435 ;
      RECT 374.185 335.705 374.385 336.435 ;
      RECT 374.685 335.705 374.885 336.435 ;
      RECT 375.18 335.705 375.38 336.435 ;
      RECT 376.475 0.17 377.245 0.43 ;
      RECT 376.475 0.17 376.735 11.5 ;
      RECT 376.985 0.17 377.245 11.5 ;
      RECT 376 335.705 376.2 336.435 ;
      RECT 376.495 335.705 376.695 336.435 ;
      RECT 377.495 0.17 378.265 0.94 ;
      RECT 377.495 0.17 377.755 12.9 ;
      RECT 378.005 0.17 378.265 12.9 ;
      RECT 376.995 335.705 377.195 336.435 ;
      RECT 377.495 335.705 377.695 336.435 ;
      RECT 377.99 335.705 378.19 336.435 ;
      RECT 378.515 0.52 378.775 5.815 ;
      RECT 379.37 0.52 379.63 5.16 ;
      RECT 379.37 4.9 380.15 5.16 ;
      RECT 379.89 4.9 380.15 6.64 ;
      RECT 378.81 335.705 379.01 336.435 ;
      RECT 379.305 335.705 379.505 336.435 ;
      RECT 379.805 335.705 380.005 336.435 ;
      RECT 380.305 335.705 380.505 336.435 ;
      RECT 380.8 335.705 381 336.435 ;
      RECT 381.62 335.705 381.82 336.435 ;
      RECT 382.115 335.705 382.315 336.435 ;
      RECT 382.615 335.705 382.815 336.435 ;
      RECT 382.77 0.52 383.03 2.335 ;
      RECT 383.115 335.705 383.315 336.435 ;
      RECT 383.28 0.52 383.54 14.11 ;
      RECT 383.61 335.705 383.81 336.435 ;
      RECT 384.655 0.17 385.425 0.94 ;
      RECT 385.165 0.17 385.425 8.7 ;
      RECT 384.655 0.17 384.915 12.9 ;
      RECT 384.145 0.52 384.405 2.485 ;
      RECT 384.43 335.705 384.63 336.435 ;
      RECT 385.675 0.17 386.445 0.43 ;
      RECT 386.185 0.17 386.445 10.48 ;
      RECT 385.675 0.17 385.935 10.99 ;
      RECT 384.925 335.705 385.125 336.435 ;
      RECT 385.425 335.705 385.625 336.435 ;
      RECT 385.925 335.705 386.125 336.435 ;
      RECT 386.42 335.705 386.62 336.435 ;
      RECT 387.715 0.17 388.485 0.43 ;
      RECT 387.715 0.17 387.975 11.5 ;
      RECT 388.225 0.17 388.485 11.5 ;
      RECT 387.24 335.705 387.44 336.435 ;
      RECT 387.735 335.705 387.935 336.435 ;
      RECT 388.735 0.17 389.505 0.94 ;
      RECT 388.735 0.17 388.995 12.9 ;
      RECT 389.245 0.17 389.505 12.9 ;
      RECT 388.235 335.705 388.435 336.435 ;
      RECT 388.735 335.705 388.935 336.435 ;
      RECT 389.23 335.705 389.43 336.435 ;
      RECT 389.755 0.52 390.015 5.815 ;
      RECT 390.61 0.52 390.87 5.16 ;
      RECT 390.61 4.9 391.39 5.16 ;
      RECT 391.13 4.9 391.39 6.64 ;
      RECT 390.05 335.705 390.25 336.435 ;
      RECT 390.545 335.705 390.745 336.435 ;
      RECT 391.045 335.705 391.245 336.435 ;
      RECT 391.545 335.705 391.745 336.435 ;
      RECT 392.04 335.705 392.24 336.435 ;
      RECT 392.86 335.705 393.06 336.435 ;
      RECT 393.355 335.705 393.555 336.435 ;
      RECT 393.855 335.705 394.055 336.435 ;
      RECT 394.01 0.52 394.27 2.335 ;
      RECT 394.355 335.705 394.555 336.435 ;
      RECT 394.52 0.52 394.78 14.11 ;
      RECT 394.85 335.705 395.05 336.435 ;
      RECT 395.895 0.17 396.665 0.94 ;
      RECT 396.405 0.17 396.665 8.7 ;
      RECT 395.895 0.17 396.155 12.9 ;
      RECT 395.385 0.52 395.645 2.485 ;
      RECT 395.67 335.705 395.87 336.435 ;
      RECT 396.915 0.17 397.685 0.43 ;
      RECT 397.425 0.17 397.685 10.48 ;
      RECT 396.915 0.17 397.175 10.99 ;
      RECT 396.165 335.705 396.365 336.435 ;
      RECT 396.665 335.705 396.865 336.435 ;
      RECT 397.165 335.705 397.365 336.435 ;
      RECT 397.66 335.705 397.86 336.435 ;
      RECT 398.955 0.17 399.725 0.43 ;
      RECT 398.955 0.17 399.215 11.5 ;
      RECT 399.465 0.17 399.725 11.5 ;
      RECT 398.48 335.705 398.68 336.435 ;
      RECT 398.975 335.705 399.175 336.435 ;
      RECT 399.975 0.17 400.745 0.94 ;
      RECT 399.975 0.17 400.235 12.9 ;
      RECT 400.485 0.17 400.745 12.9 ;
      RECT 399.475 335.705 399.675 336.435 ;
      RECT 399.975 335.705 400.175 336.435 ;
      RECT 400.47 335.705 400.67 336.435 ;
      RECT 400.995 0.52 401.255 5.815 ;
      RECT 401.85 0.52 402.11 5.16 ;
      RECT 401.85 4.9 402.63 5.16 ;
      RECT 402.37 4.9 402.63 6.64 ;
      RECT 401.29 335.705 401.49 336.435 ;
      RECT 401.785 335.705 401.985 336.435 ;
      RECT 402.285 335.705 402.485 336.435 ;
      RECT 402.785 335.705 402.985 336.435 ;
      RECT 403.28 335.705 403.48 336.435 ;
      RECT 404.1 335.705 404.3 336.435 ;
      RECT 404.595 335.705 404.795 336.435 ;
      RECT 405.095 335.705 405.295 336.435 ;
      RECT 405.25 0.52 405.51 2.335 ;
      RECT 405.595 335.705 405.795 336.435 ;
      RECT 405.76 0.52 406.02 14.11 ;
      RECT 406.09 335.705 406.29 336.435 ;
      RECT 407.135 0.17 407.905 0.94 ;
      RECT 407.645 0.17 407.905 8.7 ;
      RECT 407.135 0.17 407.395 12.9 ;
      RECT 406.625 0.52 406.885 2.485 ;
      RECT 406.91 335.705 407.11 336.435 ;
      RECT 408.155 0.17 408.925 0.43 ;
      RECT 408.665 0.17 408.925 10.48 ;
      RECT 408.155 0.17 408.415 10.99 ;
      RECT 407.405 335.705 407.605 336.435 ;
      RECT 407.905 335.705 408.105 336.435 ;
      RECT 408.405 335.705 408.605 336.435 ;
      RECT 408.9 335.705 409.1 336.435 ;
      RECT 410.195 0.17 410.965 0.43 ;
      RECT 410.195 0.17 410.455 11.5 ;
      RECT 410.705 0.17 410.965 11.5 ;
      RECT 409.72 335.705 409.92 336.435 ;
      RECT 410.215 335.705 410.415 336.435 ;
      RECT 411.215 0.17 411.985 0.94 ;
      RECT 411.215 0.17 411.475 12.9 ;
      RECT 411.725 0.17 411.985 12.9 ;
      RECT 410.715 335.705 410.915 336.435 ;
      RECT 411.215 335.705 411.415 336.435 ;
      RECT 411.71 335.705 411.91 336.435 ;
      RECT 412.235 0.52 412.495 5.815 ;
      RECT 413.09 0.52 413.35 5.16 ;
      RECT 413.09 4.9 413.87 5.16 ;
      RECT 413.61 4.9 413.87 6.64 ;
      RECT 412.53 335.705 412.73 336.435 ;
      RECT 413.025 335.705 413.225 336.435 ;
      RECT 413.525 335.705 413.725 336.435 ;
      RECT 414.025 335.705 414.225 336.435 ;
      RECT 414.52 335.705 414.72 336.435 ;
      RECT 415.34 335.705 415.54 336.435 ;
      RECT 416.335 45.465 416.535 336.435 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 272.265 0 277.095 336.46 ;
      RECT 283.505 0 288.335 336.46 ;
      RECT 294.745 0 299.575 336.46 ;
      RECT 305.985 0 310.815 336.46 ;
      RECT 317.225 0 322.055 336.46 ;
      RECT 328.465 0 333.295 336.46 ;
      RECT 339.705 0 344.535 336.46 ;
      RECT 350.945 0 355.775 336.46 ;
      RECT 362.185 0 367.015 336.46 ;
      RECT 373.425 0 378.255 336.46 ;
      RECT 384.665 0 389.495 336.46 ;
      RECT 395.905 0 400.735 336.46 ;
      RECT 407.145 0 411.975 336.46 ;
      RECT 201.98 0 202.22 336.46 ;
      RECT 203.51 0 203.75 336.46 ;
      RECT 206.57 0 206.81 336.46 ;
      RECT 208.1 0 208.34 336.46 ;
      RECT 218.3 0 222.11 336.46 ;
      RECT 223.4 0 224.15 336.46 ;
      RECT 0 0 3.03 336.46 ;
      RECT 4.655 0.17 9.505 336.46 ;
      RECT 11.65 0 14.27 336.46 ;
      RECT 15.895 0.17 20.745 336.46 ;
      RECT 22.89 0 25.51 336.46 ;
      RECT 27.135 0.17 31.985 336.46 ;
      RECT 34.13 0 36.75 336.46 ;
      RECT 38.375 0.17 43.225 336.46 ;
      RECT 45.37 0 47.99 336.46 ;
      RECT 49.615 0.17 54.465 336.46 ;
      RECT 56.61 0 59.23 336.46 ;
      RECT 60.855 0.17 65.705 336.46 ;
      RECT 67.85 0 70.47 336.46 ;
      RECT 72.095 0.17 76.945 336.46 ;
      RECT 79.09 0 81.71 336.46 ;
      RECT 83.335 0.17 88.185 336.46 ;
      RECT 90.33 0 92.95 336.46 ;
      RECT 94.575 0.17 99.425 336.46 ;
      RECT 101.57 0 104.19 336.46 ;
      RECT 105.815 0.17 110.665 336.46 ;
      RECT 112.81 0 115.43 336.46 ;
      RECT 117.055 0.17 121.905 336.46 ;
      RECT 124.05 0 126.67 336.46 ;
      RECT 128.295 0.17 133.145 336.46 ;
      RECT 135.29 0 137.91 336.46 ;
      RECT 139.535 0.17 144.385 336.46 ;
      RECT 146.53 0 149.15 336.46 ;
      RECT 150.775 0.17 155.625 336.46 ;
      RECT 157.77 0 160.39 336.46 ;
      RECT 162.015 0.17 166.865 336.46 ;
      RECT 169.01 0 171.63 336.46 ;
      RECT 173.255 0.17 178.105 336.46 ;
      RECT 180.25 0 192.03 336.46 ;
      RECT 194.32 0.17 200.7 336.46 ;
      RECT 201.97 0.3 202.23 336.46 ;
      RECT 203.5 0.3 203.76 336.46 ;
      RECT 206.56 0.3 206.82 336.46 ;
      RECT 208.09 0.3 208.35 336.46 ;
      RECT 209.63 0.17 210.9 336.46 ;
      RECT 209.62 0.3 210.9 336.46 ;
      RECT 215.23 0.17 217.02 336.46 ;
      RECT 218.29 0.3 222.12 336.46 ;
      RECT 223.39 0.3 224.16 336.46 ;
      RECT 224.93 0 236.39 336.46 ;
      RECT 224.92 0.17 236.39 336.46 ;
      RECT 238.535 0.17 243.385 336.46 ;
      RECT 245.01 0 247.63 336.46 ;
      RECT 249.775 0.17 254.625 336.46 ;
      RECT 256.25 0 258.87 336.46 ;
      RECT 261.015 0.17 265.865 336.46 ;
      RECT 267.49 0 270.11 336.46 ;
      RECT 272.255 0.17 277.105 336.46 ;
      RECT 278.73 0 281.35 336.46 ;
      RECT 283.495 0.17 288.345 336.46 ;
      RECT 289.97 0 292.59 336.46 ;
      RECT 294.735 0.17 299.585 336.46 ;
      RECT 301.21 0 303.83 336.46 ;
      RECT 305.975 0.17 310.825 336.46 ;
      RECT 312.45 0 315.07 336.46 ;
      RECT 317.215 0.17 322.065 336.46 ;
      RECT 323.69 0 326.31 336.46 ;
      RECT 328.455 0.17 333.305 336.46 ;
      RECT 334.93 0 337.55 336.46 ;
      RECT 339.695 0.17 344.545 336.46 ;
      RECT 346.17 0 348.79 336.46 ;
      RECT 350.935 0.17 355.785 336.46 ;
      RECT 357.41 0 360.03 336.46 ;
      RECT 362.175 0.17 367.025 336.46 ;
      RECT 368.65 0 371.27 336.46 ;
      RECT 373.415 0.17 378.265 336.46 ;
      RECT 379.89 0 382.51 336.46 ;
      RECT 384.655 0.17 389.505 336.46 ;
      RECT 391.13 0 393.75 336.46 ;
      RECT 395.895 0.17 400.745 336.46 ;
      RECT 402.37 0 404.99 336.46 ;
      RECT 407.135 0.17 411.985 336.46 ;
      RECT 413.61 0 416.64 336.46 ;
      RECT 0 0.52 416.64 336.46 ;
      RECT 4.665 0 9.495 336.46 ;
      RECT 15.905 0 20.735 336.46 ;
      RECT 27.145 0 31.975 336.46 ;
      RECT 38.385 0 43.215 336.46 ;
      RECT 49.625 0 54.455 336.46 ;
      RECT 60.865 0 65.695 336.46 ;
      RECT 72.105 0 76.935 336.46 ;
      RECT 83.345 0 88.175 336.46 ;
      RECT 94.585 0 99.415 336.46 ;
      RECT 105.825 0 110.655 336.46 ;
      RECT 117.065 0 121.895 336.46 ;
      RECT 128.305 0 133.135 336.46 ;
      RECT 139.545 0 144.375 336.46 ;
      RECT 150.785 0 155.615 336.46 ;
      RECT 162.025 0 166.855 336.46 ;
      RECT 173.265 0 178.095 336.46 ;
      RECT 194.32 0 200.69 336.46 ;
      RECT 209.63 0 210.89 336.46 ;
      RECT 215.23 0 217.01 336.46 ;
      RECT 238.545 0 243.375 336.46 ;
      RECT 249.785 0 254.615 336.46 ;
      RECT 261.025 0 265.855 336.46 ;
    LAYER Metal3 ;
      RECT 0 0 416.64 336.46 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 39.085 9.62 45.205 ;
      RECT 0 0 4 336.46 ;
      RECT 7.33 0 9.62 336.46 ;
      RECT 12.95 39.085 20.86 45.205 ;
      RECT 12.95 0 15.24 336.46 ;
      RECT 18.57 0 20.86 336.46 ;
      RECT 24.19 39.085 32.1 45.205 ;
      RECT 24.19 0 26.48 336.46 ;
      RECT 29.81 0 32.1 336.46 ;
      RECT 35.43 39.085 43.34 45.205 ;
      RECT 35.43 0 37.72 336.46 ;
      RECT 41.05 0 43.34 336.46 ;
      RECT 46.67 39.085 54.58 45.205 ;
      RECT 46.67 0 48.96 336.46 ;
      RECT 52.29 0 54.58 336.46 ;
      RECT 57.91 39.085 65.82 45.205 ;
      RECT 57.91 0 60.2 336.46 ;
      RECT 63.53 0 65.82 336.46 ;
      RECT 69.15 39.085 77.06 45.205 ;
      RECT 69.15 0 71.44 336.46 ;
      RECT 74.77 0 77.06 336.46 ;
      RECT 80.39 39.085 88.3 45.205 ;
      RECT 80.39 0 82.68 336.46 ;
      RECT 86.01 0 88.3 336.46 ;
      RECT 91.63 39.085 99.54 45.205 ;
      RECT 91.63 0 93.92 336.46 ;
      RECT 97.25 0 99.54 336.46 ;
      RECT 102.87 39.085 110.78 45.205 ;
      RECT 102.87 0 105.16 336.46 ;
      RECT 108.49 0 110.78 336.46 ;
      RECT 114.11 39.085 122.02 45.205 ;
      RECT 114.11 0 116.4 336.46 ;
      RECT 119.73 0 122.02 336.46 ;
      RECT 125.35 39.085 133.26 45.205 ;
      RECT 125.35 0 127.64 336.46 ;
      RECT 130.97 0 133.26 336.46 ;
      RECT 136.59 39.085 144.5 45.205 ;
      RECT 136.59 0 138.88 336.46 ;
      RECT 142.21 0 144.5 336.46 ;
      RECT 147.83 39.085 155.74 45.205 ;
      RECT 147.83 0 150.12 336.46 ;
      RECT 153.45 0 155.74 336.46 ;
      RECT 159.07 39.085 166.98 45.205 ;
      RECT 159.07 0 161.36 336.46 ;
      RECT 164.69 0 166.98 336.46 ;
      RECT 170.31 39.085 178.22 45.205 ;
      RECT 170.31 0 172.6 336.46 ;
      RECT 175.93 0 178.22 336.46 ;
      RECT 181.55 0 188.63 336.46 ;
      RECT 191.96 0 193.78 336.46 ;
      RECT 197.11 0 198.93 336.46 ;
      RECT 202.26 0 204.08 336.46 ;
      RECT 207.41 0 209.23 336.46 ;
      RECT 212.56 0 214.38 336.46 ;
      RECT 238.42 39.085 246.33 45.205 ;
      RECT 238.42 0 240.71 336.46 ;
      RECT 244.04 0 246.33 336.46 ;
      RECT 249.66 39.085 257.57 45.205 ;
      RECT 249.66 0 251.95 336.46 ;
      RECT 255.28 0 257.57 336.46 ;
      RECT 260.9 39.085 268.81 45.205 ;
      RECT 260.9 0 263.19 336.46 ;
      RECT 266.52 0 268.81 336.46 ;
      RECT 272.14 39.085 280.05 45.205 ;
      RECT 272.14 0 274.43 336.46 ;
      RECT 277.76 0 280.05 336.46 ;
      RECT 283.38 39.085 291.29 45.205 ;
      RECT 283.38 0 285.67 336.46 ;
      RECT 289 0 291.29 336.46 ;
      RECT 294.62 39.085 302.53 45.205 ;
      RECT 294.62 0 296.91 336.46 ;
      RECT 300.24 0 302.53 336.46 ;
      RECT 305.86 39.085 313.77 45.205 ;
      RECT 305.86 0 308.15 336.46 ;
      RECT 311.48 0 313.77 336.46 ;
      RECT 317.1 39.085 325.01 45.205 ;
      RECT 317.1 0 319.39 336.46 ;
      RECT 322.72 0 325.01 336.46 ;
      RECT 328.34 39.085 336.25 45.205 ;
      RECT 328.34 0 330.63 336.46 ;
      RECT 333.96 0 336.25 336.46 ;
      RECT 339.58 39.085 347.49 45.205 ;
      RECT 339.58 0 341.87 336.46 ;
      RECT 345.2 0 347.49 336.46 ;
      RECT 350.82 39.085 358.73 45.205 ;
      RECT 350.82 0 353.11 336.46 ;
      RECT 356.44 0 358.73 336.46 ;
      RECT 362.06 39.085 369.97 45.205 ;
      RECT 362.06 0 364.35 336.46 ;
      RECT 367.68 0 369.97 336.46 ;
      RECT 373.3 39.085 381.21 45.205 ;
      RECT 373.3 0 375.59 336.46 ;
      RECT 378.92 0 381.21 336.46 ;
      RECT 384.54 39.085 392.45 45.205 ;
      RECT 384.54 0 386.83 336.46 ;
      RECT 390.16 0 392.45 336.46 ;
      RECT 395.78 39.085 403.69 45.205 ;
      RECT 395.78 0 398.07 336.46 ;
      RECT 401.4 0 403.69 336.46 ;
      RECT 407.02 39.085 416.64 45.205 ;
      RECT 407.02 0 409.31 336.46 ;
      RECT 412.64 0 416.64 336.46 ;
      RECT 217.71 0 219.53 336.46 ;
      RECT 222.86 0 224.68 336.46 ;
      RECT 228.01 0 235.09 336.46 ;
  END
END RM_IHPSG13_1P_1024x32_c2_bm_bist

END LIBRARY
