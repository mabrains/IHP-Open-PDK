# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 16:22:45 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_256x8_c3_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_256x8_c3_bm_bist 0 0 ;
  SIZE 236.8 BY 74.1 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.09 0 155.35 0.26 ;
    END
  END A_DIN[4]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.45 0 81.71 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.56 0 153.82 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.98 0 83.24 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 158.97 0 159.23 0.26 ;
    END
  END A_BM[4]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.57 0 77.83 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.5 0 160.76 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.04 0 76.3 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 159.835 0 160.095 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.705 0 76.965 0.26 ;
    END
  END A_DOUT[3]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 224.11 0 226.92 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.87 0 215.68 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 201.63 0 204.44 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.39 0 193.2 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.15 0 181.96 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.91 0 170.72 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.67 0 159.48 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.43 0 148.24 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.02 0 137.83 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.72 0 127.53 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.27 0 112.08 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 98.97 0 101.78 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 74.1 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 0 232.54 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 0 221.3 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 0 210.06 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 0 198.82 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 0 187.58 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 0 176.34 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 0 165.1 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 0 153.86 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.87 0 132.68 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.57 0 122.38 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 114.42 0 117.23 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 104.12 0 106.93 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 30.425 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 229.73 37.065 232.54 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.49 37.065 221.3 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 207.25 37.065 210.06 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 196.01 37.065 198.82 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.77 37.065 187.58 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 173.53 37.065 176.34 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 162.29 37.065 165.1 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.05 37.065 153.86 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 37.065 85.75 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 37.065 74.51 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 37.065 63.27 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 37.065 52.03 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 37.065 40.79 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 37.065 29.55 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 37.065 18.31 74.1 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 37.065 7.07 74.1 ;
    END
  END VDDARRAY!
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 177.57 0 177.83 0.26 ;
    END
  END A_DIN[5]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 58.97 0 59.23 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.04 0 176.3 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.5 0 60.76 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.45 0 181.71 0.26 ;
    END
  END A_BM[5]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.09 0 55.35 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.98 0 183.24 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.56 0 53.82 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.315 0 182.575 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.225 0 54.485 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.05 0 200.31 0.26 ;
    END
  END A_DIN[6]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.49 0 36.75 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 198.52 0 198.78 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.02 0 38.28 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.93 0 204.19 0.26 ;
    END
  END A_BM[6]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.61 0 32.87 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.46 0 205.72 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.08 0 31.34 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.795 0 205.055 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.745 0 32.005 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 222.53 0 222.79 0.26 ;
    END
  END A_DIN[7]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.01 0 14.27 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221 0 221.26 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.54 0 15.8 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 226.41 0 226.67 0.26 ;
    END
  END A_BM[7]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.13 0 10.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.94 0 228.2 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 8.6 0 8.86 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.275 0 227.535 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.265 0 9.525 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7171 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 34.349515 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.6 0 114.86 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5127 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 38.31068 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.19 0 119.45 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.59 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 28.783172 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.09 0 114.35 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3856 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 32.744337 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 118.68 0 118.94 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4519 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 33.029126 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.81 0 100.07 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1867 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 31.708738 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.34 0 101.6 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.25 0 122.51 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 122.76 0 123.02 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.23 0 121.49 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 121.74 0 122 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0139 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.763754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.8 0 125.06 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7487 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.443366 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.29 0 124.55 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7429 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 59.372168 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.78 0 124.04 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4777 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 58.05178 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.27 0 123.53 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.36 0 102.62 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4931 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.191934 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.87 0 103.13 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8707 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.220065 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.56 0 112.82 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81105 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.923077 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.13 0 116.39 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.62 0 115.88 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8407 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.09186 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.07 0 113.33 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.874 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 12.046332 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.49 0 134.75 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 72.69295 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.01 LAYER Metal3 ;
      ANTENNAMAXAREACAR 1.686364 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.344457 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.11 0 115.37 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9799 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 11.079661 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.03 0 111.29 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9279 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.820762 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.66 0 117.92 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7211 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.812298 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.15 0 117.41 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7137 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.775454 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.54 0 111.8 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 236.8 74.1 ;
    LAYER Metal2 ;
      RECT 0.105 37.065 0.305 74.075 ;
      RECT 1.1 73.345 1.3 74.075 ;
      RECT 1.92 73.345 2.12 74.075 ;
      RECT 2.415 73.345 2.615 74.075 ;
      RECT 2.915 73.345 3.115 74.075 ;
      RECT 3.415 73.345 3.615 74.075 ;
      RECT 3.91 73.345 4.11 74.075 ;
      RECT 4.73 73.345 4.93 74.075 ;
      RECT 5.225 73.345 5.425 74.075 ;
      RECT 5.725 73.345 5.925 74.075 ;
      RECT 7.225 0.17 7.995 0.43 ;
      RECT 7.225 0.17 7.485 11.38 ;
      RECT 7.735 0.17 7.995 17.1 ;
      RECT 6.225 73.345 6.425 74.075 ;
      RECT 6.72 73.345 6.92 74.075 ;
      RECT 7.54 73.345 7.74 74.075 ;
      RECT 8.035 73.345 8.235 74.075 ;
      RECT 8.535 73.345 8.735 74.075 ;
      RECT 8.6 0.52 8.86 2.255 ;
      RECT 9.035 73.345 9.235 74.075 ;
      RECT 9.265 0.52 9.525 8.085 ;
      RECT 9.53 73.345 9.73 74.075 ;
      RECT 10.13 0.52 10.39 1.5 ;
      RECT 10.35 73.345 10.55 74.075 ;
      RECT 10.845 73.345 11.045 74.075 ;
      RECT 11.345 73.345 11.545 74.075 ;
      RECT 11.845 73.345 12.045 74.075 ;
      RECT 12.34 73.345 12.54 74.075 ;
      RECT 13.16 73.345 13.36 74.075 ;
      RECT 13.655 73.345 13.855 74.075 ;
      RECT 14.01 0.52 14.27 2.255 ;
      RECT 14.155 73.345 14.355 74.075 ;
      RECT 14.655 73.345 14.855 74.075 ;
      RECT 15.15 73.345 15.35 74.075 ;
      RECT 16.255 0.8 17.025 1.57 ;
      RECT 16.255 0.3 16.515 13.03 ;
      RECT 16.765 0.3 17.025 13.03 ;
      RECT 15.54 0.52 15.8 2.255 ;
      RECT 15.97 73.345 16.17 74.075 ;
      RECT 16.465 73.345 16.665 74.075 ;
      RECT 16.965 73.345 17.165 74.075 ;
      RECT 17.465 73.345 17.665 74.075 ;
      RECT 17.96 73.345 18.16 74.075 ;
      RECT 18.78 73.345 18.98 74.075 ;
      RECT 19.975 0.17 20.745 0.43 ;
      RECT 19.975 0.17 20.235 13.055 ;
      RECT 20.485 0.17 20.745 13.055 ;
      RECT 19.275 73.345 19.475 74.075 ;
      RECT 19.775 73.345 19.975 74.075 ;
      RECT 20.275 73.345 20.475 74.075 ;
      RECT 20.77 73.345 20.97 74.075 ;
      RECT 21.59 73.345 21.79 74.075 ;
      RECT 22.085 73.345 22.285 74.075 ;
      RECT 22.585 73.345 22.785 74.075 ;
      RECT 23.085 73.345 23.285 74.075 ;
      RECT 23.58 73.345 23.78 74.075 ;
      RECT 24.4 73.345 24.6 74.075 ;
      RECT 24.895 73.345 25.095 74.075 ;
      RECT 25.395 73.345 25.595 74.075 ;
      RECT 25.895 73.345 26.095 74.075 ;
      RECT 26.39 73.345 26.59 74.075 ;
      RECT 27.21 73.345 27.41 74.075 ;
      RECT 27.705 73.345 27.905 74.075 ;
      RECT 28.205 73.345 28.405 74.075 ;
      RECT 29.705 0.17 30.475 0.43 ;
      RECT 29.705 0.17 29.965 11.38 ;
      RECT 30.215 0.17 30.475 17.1 ;
      RECT 28.705 73.345 28.905 74.075 ;
      RECT 29.2 73.345 29.4 74.075 ;
      RECT 30.02 73.345 30.22 74.075 ;
      RECT 30.515 73.345 30.715 74.075 ;
      RECT 31.015 73.345 31.215 74.075 ;
      RECT 31.08 0.52 31.34 2.255 ;
      RECT 31.515 73.345 31.715 74.075 ;
      RECT 31.745 0.52 32.005 8.085 ;
      RECT 32.01 73.345 32.21 74.075 ;
      RECT 32.61 0.52 32.87 1.5 ;
      RECT 32.83 73.345 33.03 74.075 ;
      RECT 33.325 73.345 33.525 74.075 ;
      RECT 33.825 73.345 34.025 74.075 ;
      RECT 34.325 73.345 34.525 74.075 ;
      RECT 34.82 73.345 35.02 74.075 ;
      RECT 35.64 73.345 35.84 74.075 ;
      RECT 36.135 73.345 36.335 74.075 ;
      RECT 36.49 0.52 36.75 2.255 ;
      RECT 36.635 73.345 36.835 74.075 ;
      RECT 37.135 73.345 37.335 74.075 ;
      RECT 37.63 73.345 37.83 74.075 ;
      RECT 38.735 0.8 39.505 1.57 ;
      RECT 38.735 0.3 38.995 13.03 ;
      RECT 39.245 0.3 39.505 13.03 ;
      RECT 38.02 0.52 38.28 2.255 ;
      RECT 38.45 73.345 38.65 74.075 ;
      RECT 38.945 73.345 39.145 74.075 ;
      RECT 39.445 73.345 39.645 74.075 ;
      RECT 39.945 73.345 40.145 74.075 ;
      RECT 40.44 73.345 40.64 74.075 ;
      RECT 41.26 73.345 41.46 74.075 ;
      RECT 42.455 0.17 43.225 0.43 ;
      RECT 42.455 0.17 42.715 13.055 ;
      RECT 42.965 0.17 43.225 13.055 ;
      RECT 41.755 73.345 41.955 74.075 ;
      RECT 42.255 73.345 42.455 74.075 ;
      RECT 42.755 73.345 42.955 74.075 ;
      RECT 43.25 73.345 43.45 74.075 ;
      RECT 44.07 73.345 44.27 74.075 ;
      RECT 44.565 73.345 44.765 74.075 ;
      RECT 45.065 73.345 45.265 74.075 ;
      RECT 45.565 73.345 45.765 74.075 ;
      RECT 46.06 73.345 46.26 74.075 ;
      RECT 46.88 73.345 47.08 74.075 ;
      RECT 47.375 73.345 47.575 74.075 ;
      RECT 47.875 73.345 48.075 74.075 ;
      RECT 48.375 73.345 48.575 74.075 ;
      RECT 48.87 73.345 49.07 74.075 ;
      RECT 49.69 73.345 49.89 74.075 ;
      RECT 50.185 73.345 50.385 74.075 ;
      RECT 50.685 73.345 50.885 74.075 ;
      RECT 52.185 0.17 52.955 0.43 ;
      RECT 52.185 0.17 52.445 11.38 ;
      RECT 52.695 0.17 52.955 17.1 ;
      RECT 51.185 73.345 51.385 74.075 ;
      RECT 51.68 73.345 51.88 74.075 ;
      RECT 52.5 73.345 52.7 74.075 ;
      RECT 52.995 73.345 53.195 74.075 ;
      RECT 53.495 73.345 53.695 74.075 ;
      RECT 53.56 0.52 53.82 2.255 ;
      RECT 53.995 73.345 54.195 74.075 ;
      RECT 54.225 0.52 54.485 8.085 ;
      RECT 54.49 73.345 54.69 74.075 ;
      RECT 55.09 0.52 55.35 1.5 ;
      RECT 55.31 73.345 55.51 74.075 ;
      RECT 55.805 73.345 56.005 74.075 ;
      RECT 56.305 73.345 56.505 74.075 ;
      RECT 56.805 73.345 57.005 74.075 ;
      RECT 57.3 73.345 57.5 74.075 ;
      RECT 58.12 73.345 58.32 74.075 ;
      RECT 58.615 73.345 58.815 74.075 ;
      RECT 58.97 0.52 59.23 2.255 ;
      RECT 59.115 73.345 59.315 74.075 ;
      RECT 59.615 73.345 59.815 74.075 ;
      RECT 60.11 73.345 60.31 74.075 ;
      RECT 61.215 0.8 61.985 1.57 ;
      RECT 61.215 0.3 61.475 13.03 ;
      RECT 61.725 0.3 61.985 13.03 ;
      RECT 60.5 0.52 60.76 2.255 ;
      RECT 60.93 73.345 61.13 74.075 ;
      RECT 61.425 73.345 61.625 74.075 ;
      RECT 61.925 73.345 62.125 74.075 ;
      RECT 62.425 73.345 62.625 74.075 ;
      RECT 62.92 73.345 63.12 74.075 ;
      RECT 63.74 73.345 63.94 74.075 ;
      RECT 64.935 0.17 65.705 0.43 ;
      RECT 64.935 0.17 65.195 13.055 ;
      RECT 65.445 0.17 65.705 13.055 ;
      RECT 64.235 73.345 64.435 74.075 ;
      RECT 64.735 73.345 64.935 74.075 ;
      RECT 65.235 73.345 65.435 74.075 ;
      RECT 65.73 73.345 65.93 74.075 ;
      RECT 66.55 73.345 66.75 74.075 ;
      RECT 67.045 73.345 67.245 74.075 ;
      RECT 67.545 73.345 67.745 74.075 ;
      RECT 68.045 73.345 68.245 74.075 ;
      RECT 68.54 73.345 68.74 74.075 ;
      RECT 69.36 73.345 69.56 74.075 ;
      RECT 69.855 73.345 70.055 74.075 ;
      RECT 70.355 73.345 70.555 74.075 ;
      RECT 70.855 73.345 71.055 74.075 ;
      RECT 71.35 73.345 71.55 74.075 ;
      RECT 72.17 73.345 72.37 74.075 ;
      RECT 72.665 73.345 72.865 74.075 ;
      RECT 73.165 73.345 73.365 74.075 ;
      RECT 74.665 0.17 75.435 0.43 ;
      RECT 74.665 0.17 74.925 11.38 ;
      RECT 75.175 0.17 75.435 17.1 ;
      RECT 73.665 73.345 73.865 74.075 ;
      RECT 74.16 73.345 74.36 74.075 ;
      RECT 74.98 73.345 75.18 74.075 ;
      RECT 75.475 73.345 75.675 74.075 ;
      RECT 75.975 73.345 76.175 74.075 ;
      RECT 76.04 0.52 76.3 2.255 ;
      RECT 76.475 73.345 76.675 74.075 ;
      RECT 76.705 0.52 76.965 8.085 ;
      RECT 76.97 73.345 77.17 74.075 ;
      RECT 77.57 0.52 77.83 1.5 ;
      RECT 77.79 73.345 77.99 74.075 ;
      RECT 78.285 73.345 78.485 74.075 ;
      RECT 78.785 73.345 78.985 74.075 ;
      RECT 79.285 73.345 79.485 74.075 ;
      RECT 79.78 73.345 79.98 74.075 ;
      RECT 80.6 73.345 80.8 74.075 ;
      RECT 81.095 73.345 81.295 74.075 ;
      RECT 81.45 0.52 81.71 2.255 ;
      RECT 81.595 73.345 81.795 74.075 ;
      RECT 82.095 73.345 82.295 74.075 ;
      RECT 82.59 73.345 82.79 74.075 ;
      RECT 83.695 0.8 84.465 1.57 ;
      RECT 83.695 0.3 83.955 13.03 ;
      RECT 84.205 0.3 84.465 13.03 ;
      RECT 82.98 0.52 83.24 2.255 ;
      RECT 83.41 73.345 83.61 74.075 ;
      RECT 83.905 73.345 84.105 74.075 ;
      RECT 84.405 73.345 84.605 74.075 ;
      RECT 84.905 73.345 85.105 74.075 ;
      RECT 85.4 73.345 85.6 74.075 ;
      RECT 86.22 73.345 86.42 74.075 ;
      RECT 87.415 0.17 88.185 0.43 ;
      RECT 87.415 0.17 87.675 13.055 ;
      RECT 87.925 0.17 88.185 13.055 ;
      RECT 86.715 73.345 86.915 74.075 ;
      RECT 87.215 73.345 87.415 74.075 ;
      RECT 87.715 73.345 87.915 74.075 ;
      RECT 88.21 73.345 88.41 74.075 ;
      RECT 89.03 73.345 89.23 74.075 ;
      RECT 89.525 73.345 89.725 74.075 ;
      RECT 90.025 73.345 90.225 74.075 ;
      RECT 90.525 73.345 90.725 74.075 ;
      RECT 96.595 0.17 97.365 0.43 ;
      RECT 96.595 0.17 96.855 36.945 ;
      RECT 97.105 0.17 97.365 36.945 ;
      RECT 91.02 73.345 91.22 74.075 ;
      RECT 91.84 73.345 92.04 74.075 ;
      RECT 99.3 0 99.56 4.94 ;
      RECT 99.3 4.68 100.07 4.94 ;
      RECT 99.81 4.68 100.07 12.9 ;
      RECT 99.81 0.52 100.07 1.78 ;
      RECT 99.81 1.52 100.58 1.78 ;
      RECT 100.32 1.52 100.58 12.9 ;
      RECT 92.835 73.345 93.035 74.075 ;
      RECT 100.32 0.59 101.09 1.27 ;
      RECT 100.83 0.59 101.09 7.965 ;
      RECT 97.615 0.3 97.875 37.365 ;
      RECT 98.125 0.3 98.385 37.365 ;
      RECT 101.34 0.52 101.6 12.9 ;
      RECT 101.85 0 102.11 12.9 ;
      RECT 102.36 0.52 102.62 12.9 ;
      RECT 102.87 0.52 103.13 12.9 ;
      RECT 103.38 0 103.64 12.9 ;
      RECT 106.44 0.17 107.21 0.43 ;
      RECT 106.44 0.17 106.7 2.085 ;
      RECT 106.95 0.17 107.21 9 ;
      RECT 103.89 0 104.15 12.9 ;
      RECT 104.4 0 104.66 8.565 ;
      RECT 104.91 0 105.17 8.055 ;
      RECT 111.03 0.52 111.29 6.59 ;
      RECT 112.56 0.52 112.82 6.305 ;
      RECT 112.56 6.045 113.53 6.305 ;
      RECT 111.54 0.52 111.8 2.23 ;
      RECT 113.07 0.52 113.33 2.955 ;
      RECT 114.09 0.52 114.35 12.9 ;
      RECT 114.6 0.52 114.86 12.9 ;
      RECT 116.13 0.52 116.39 6.29 ;
      RECT 115.62 6.045 116.39 6.29 ;
      RECT 115.11 0.52 115.37 6.745 ;
      RECT 117.66 0.52 117.92 6.59 ;
      RECT 117.015 6.33 117.92 6.59 ;
      RECT 115.62 0.52 115.88 2.955 ;
      RECT 117.15 0.52 117.41 2.67 ;
      RECT 118.68 0.52 118.94 12.9 ;
      RECT 119.19 0.52 119.45 12.9 ;
      RECT 120.72 0.575 120.98 7.965 ;
      RECT 121.23 0.52 121.49 12.9 ;
      RECT 121.74 0.52 122 12.9 ;
      RECT 122.25 0.52 122.51 12.9 ;
      RECT 122.76 0.52 123.02 12.9 ;
      RECT 123.27 0.52 123.53 12.9 ;
      RECT 123.78 0.52 124.04 12.9 ;
      RECT 124.29 0.52 124.55 12.9 ;
      RECT 124.8 0.52 125.06 12.9 ;
      RECT 125.31 0 125.57 12.9 ;
      RECT 125.82 0 126.08 12.9 ;
      RECT 127.35 0 127.61 12.9 ;
      RECT 127.86 0 128.12 12.9 ;
      RECT 135 0.17 135.77 0.43 ;
      RECT 135 0.17 135.26 13.845 ;
      RECT 135.51 0.17 135.77 13.845 ;
      RECT 137.04 0.17 137.81 0.43 ;
      RECT 137.04 0.17 137.3 2.11 ;
      RECT 137.55 0.17 137.81 2.11 ;
      RECT 132.45 0 132.71 3.61 ;
      RECT 132.96 0 133.22 4.12 ;
      RECT 139.435 0.17 140.205 0.43 ;
      RECT 139.435 0.17 139.695 36.945 ;
      RECT 139.945 0.17 140.205 36.945 ;
      RECT 134.49 0.52 134.75 15.16 ;
      RECT 138.415 0.3 138.675 37.365 ;
      RECT 138.925 0.3 139.185 37.365 ;
      RECT 143.765 73.345 143.965 74.075 ;
      RECT 144.76 73.345 144.96 74.075 ;
      RECT 145.58 73.345 145.78 74.075 ;
      RECT 146.075 73.345 146.275 74.075 ;
      RECT 146.575 73.345 146.775 74.075 ;
      RECT 147.075 73.345 147.275 74.075 ;
      RECT 148.615 0.17 149.385 0.43 ;
      RECT 148.615 0.17 148.875 13.055 ;
      RECT 149.125 0.17 149.385 13.055 ;
      RECT 147.57 73.345 147.77 74.075 ;
      RECT 148.39 73.345 148.59 74.075 ;
      RECT 148.885 73.345 149.085 74.075 ;
      RECT 149.385 73.345 149.585 74.075 ;
      RECT 149.885 73.345 150.085 74.075 ;
      RECT 150.38 73.345 150.58 74.075 ;
      RECT 151.2 73.345 151.4 74.075 ;
      RECT 152.335 0.8 153.105 1.57 ;
      RECT 152.335 0.3 152.595 13.03 ;
      RECT 152.845 0.3 153.105 13.03 ;
      RECT 151.695 73.345 151.895 74.075 ;
      RECT 152.195 73.345 152.395 74.075 ;
      RECT 152.695 73.345 152.895 74.075 ;
      RECT 153.19 73.345 153.39 74.075 ;
      RECT 153.56 0.52 153.82 2.255 ;
      RECT 154.01 73.345 154.21 74.075 ;
      RECT 154.505 73.345 154.705 74.075 ;
      RECT 155.005 73.345 155.205 74.075 ;
      RECT 155.09 0.52 155.35 2.255 ;
      RECT 155.505 73.345 155.705 74.075 ;
      RECT 156 73.345 156.2 74.075 ;
      RECT 156.82 73.345 157.02 74.075 ;
      RECT 157.315 73.345 157.515 74.075 ;
      RECT 157.815 73.345 158.015 74.075 ;
      RECT 158.315 73.345 158.515 74.075 ;
      RECT 158.81 73.345 159.01 74.075 ;
      RECT 158.97 0.52 159.23 1.5 ;
      RECT 159.63 73.345 159.83 74.075 ;
      RECT 159.835 0.52 160.095 8.085 ;
      RECT 160.125 73.345 160.325 74.075 ;
      RECT 160.5 0.52 160.76 2.255 ;
      RECT 161.365 0.17 162.135 0.43 ;
      RECT 161.875 0.17 162.135 11.38 ;
      RECT 161.365 0.17 161.625 17.1 ;
      RECT 160.625 73.345 160.825 74.075 ;
      RECT 161.125 73.345 161.325 74.075 ;
      RECT 161.62 73.345 161.82 74.075 ;
      RECT 162.44 73.345 162.64 74.075 ;
      RECT 162.935 73.345 163.135 74.075 ;
      RECT 163.435 73.345 163.635 74.075 ;
      RECT 163.935 73.345 164.135 74.075 ;
      RECT 164.43 73.345 164.63 74.075 ;
      RECT 165.25 73.345 165.45 74.075 ;
      RECT 165.745 73.345 165.945 74.075 ;
      RECT 166.245 73.345 166.445 74.075 ;
      RECT 166.745 73.345 166.945 74.075 ;
      RECT 167.24 73.345 167.44 74.075 ;
      RECT 168.06 73.345 168.26 74.075 ;
      RECT 168.555 73.345 168.755 74.075 ;
      RECT 169.055 73.345 169.255 74.075 ;
      RECT 169.555 73.345 169.755 74.075 ;
      RECT 171.095 0.17 171.865 0.43 ;
      RECT 171.095 0.17 171.355 13.055 ;
      RECT 171.605 0.17 171.865 13.055 ;
      RECT 170.05 73.345 170.25 74.075 ;
      RECT 170.87 73.345 171.07 74.075 ;
      RECT 171.365 73.345 171.565 74.075 ;
      RECT 171.865 73.345 172.065 74.075 ;
      RECT 172.365 73.345 172.565 74.075 ;
      RECT 172.86 73.345 173.06 74.075 ;
      RECT 173.68 73.345 173.88 74.075 ;
      RECT 174.815 0.8 175.585 1.57 ;
      RECT 174.815 0.3 175.075 13.03 ;
      RECT 175.325 0.3 175.585 13.03 ;
      RECT 174.175 73.345 174.375 74.075 ;
      RECT 174.675 73.345 174.875 74.075 ;
      RECT 175.175 73.345 175.375 74.075 ;
      RECT 175.67 73.345 175.87 74.075 ;
      RECT 176.04 0.52 176.3 2.255 ;
      RECT 176.49 73.345 176.69 74.075 ;
      RECT 176.985 73.345 177.185 74.075 ;
      RECT 177.485 73.345 177.685 74.075 ;
      RECT 177.57 0.52 177.83 2.255 ;
      RECT 177.985 73.345 178.185 74.075 ;
      RECT 178.48 73.345 178.68 74.075 ;
      RECT 179.3 73.345 179.5 74.075 ;
      RECT 179.795 73.345 179.995 74.075 ;
      RECT 180.295 73.345 180.495 74.075 ;
      RECT 180.795 73.345 180.995 74.075 ;
      RECT 181.29 73.345 181.49 74.075 ;
      RECT 181.45 0.52 181.71 1.5 ;
      RECT 182.11 73.345 182.31 74.075 ;
      RECT 182.315 0.52 182.575 8.085 ;
      RECT 182.605 73.345 182.805 74.075 ;
      RECT 182.98 0.52 183.24 2.255 ;
      RECT 183.845 0.17 184.615 0.43 ;
      RECT 184.355 0.17 184.615 11.38 ;
      RECT 183.845 0.17 184.105 17.1 ;
      RECT 183.105 73.345 183.305 74.075 ;
      RECT 183.605 73.345 183.805 74.075 ;
      RECT 184.1 73.345 184.3 74.075 ;
      RECT 184.92 73.345 185.12 74.075 ;
      RECT 185.415 73.345 185.615 74.075 ;
      RECT 185.915 73.345 186.115 74.075 ;
      RECT 186.415 73.345 186.615 74.075 ;
      RECT 186.91 73.345 187.11 74.075 ;
      RECT 187.73 73.345 187.93 74.075 ;
      RECT 188.225 73.345 188.425 74.075 ;
      RECT 188.725 73.345 188.925 74.075 ;
      RECT 189.225 73.345 189.425 74.075 ;
      RECT 189.72 73.345 189.92 74.075 ;
      RECT 190.54 73.345 190.74 74.075 ;
      RECT 191.035 73.345 191.235 74.075 ;
      RECT 191.535 73.345 191.735 74.075 ;
      RECT 192.035 73.345 192.235 74.075 ;
      RECT 193.575 0.17 194.345 0.43 ;
      RECT 193.575 0.17 193.835 13.055 ;
      RECT 194.085 0.17 194.345 13.055 ;
      RECT 192.53 73.345 192.73 74.075 ;
      RECT 193.35 73.345 193.55 74.075 ;
      RECT 193.845 73.345 194.045 74.075 ;
      RECT 194.345 73.345 194.545 74.075 ;
      RECT 194.845 73.345 195.045 74.075 ;
      RECT 195.34 73.345 195.54 74.075 ;
      RECT 196.16 73.345 196.36 74.075 ;
      RECT 197.295 0.8 198.065 1.57 ;
      RECT 197.295 0.3 197.555 13.03 ;
      RECT 197.805 0.3 198.065 13.03 ;
      RECT 196.655 73.345 196.855 74.075 ;
      RECT 197.155 73.345 197.355 74.075 ;
      RECT 197.655 73.345 197.855 74.075 ;
      RECT 198.15 73.345 198.35 74.075 ;
      RECT 198.52 0.52 198.78 2.255 ;
      RECT 198.97 73.345 199.17 74.075 ;
      RECT 199.465 73.345 199.665 74.075 ;
      RECT 199.965 73.345 200.165 74.075 ;
      RECT 200.05 0.52 200.31 2.255 ;
      RECT 200.465 73.345 200.665 74.075 ;
      RECT 200.96 73.345 201.16 74.075 ;
      RECT 201.78 73.345 201.98 74.075 ;
      RECT 202.275 73.345 202.475 74.075 ;
      RECT 202.775 73.345 202.975 74.075 ;
      RECT 203.275 73.345 203.475 74.075 ;
      RECT 203.77 73.345 203.97 74.075 ;
      RECT 203.93 0.52 204.19 1.5 ;
      RECT 204.59 73.345 204.79 74.075 ;
      RECT 204.795 0.52 205.055 8.085 ;
      RECT 205.085 73.345 205.285 74.075 ;
      RECT 205.46 0.52 205.72 2.255 ;
      RECT 206.325 0.17 207.095 0.43 ;
      RECT 206.835 0.17 207.095 11.38 ;
      RECT 206.325 0.17 206.585 17.1 ;
      RECT 205.585 73.345 205.785 74.075 ;
      RECT 206.085 73.345 206.285 74.075 ;
      RECT 206.58 73.345 206.78 74.075 ;
      RECT 207.4 73.345 207.6 74.075 ;
      RECT 207.895 73.345 208.095 74.075 ;
      RECT 208.395 73.345 208.595 74.075 ;
      RECT 208.895 73.345 209.095 74.075 ;
      RECT 209.39 73.345 209.59 74.075 ;
      RECT 210.21 73.345 210.41 74.075 ;
      RECT 210.705 73.345 210.905 74.075 ;
      RECT 211.205 73.345 211.405 74.075 ;
      RECT 211.705 73.345 211.905 74.075 ;
      RECT 212.2 73.345 212.4 74.075 ;
      RECT 213.02 73.345 213.22 74.075 ;
      RECT 213.515 73.345 213.715 74.075 ;
      RECT 214.015 73.345 214.215 74.075 ;
      RECT 214.515 73.345 214.715 74.075 ;
      RECT 216.055 0.17 216.825 0.43 ;
      RECT 216.055 0.17 216.315 13.055 ;
      RECT 216.565 0.17 216.825 13.055 ;
      RECT 215.01 73.345 215.21 74.075 ;
      RECT 215.83 73.345 216.03 74.075 ;
      RECT 216.325 73.345 216.525 74.075 ;
      RECT 216.825 73.345 217.025 74.075 ;
      RECT 217.325 73.345 217.525 74.075 ;
      RECT 217.82 73.345 218.02 74.075 ;
      RECT 218.64 73.345 218.84 74.075 ;
      RECT 219.775 0.8 220.545 1.57 ;
      RECT 219.775 0.3 220.035 13.03 ;
      RECT 220.285 0.3 220.545 13.03 ;
      RECT 219.135 73.345 219.335 74.075 ;
      RECT 219.635 73.345 219.835 74.075 ;
      RECT 220.135 73.345 220.335 74.075 ;
      RECT 220.63 73.345 220.83 74.075 ;
      RECT 221 0.52 221.26 2.255 ;
      RECT 221.45 73.345 221.65 74.075 ;
      RECT 221.945 73.345 222.145 74.075 ;
      RECT 222.445 73.345 222.645 74.075 ;
      RECT 222.53 0.52 222.79 2.255 ;
      RECT 222.945 73.345 223.145 74.075 ;
      RECT 223.44 73.345 223.64 74.075 ;
      RECT 224.26 73.345 224.46 74.075 ;
      RECT 224.755 73.345 224.955 74.075 ;
      RECT 225.255 73.345 225.455 74.075 ;
      RECT 225.755 73.345 225.955 74.075 ;
      RECT 226.25 73.345 226.45 74.075 ;
      RECT 226.41 0.52 226.67 1.5 ;
      RECT 227.07 73.345 227.27 74.075 ;
      RECT 227.275 0.52 227.535 8.085 ;
      RECT 227.565 73.345 227.765 74.075 ;
      RECT 227.94 0.52 228.2 2.255 ;
      RECT 228.805 0.17 229.575 0.43 ;
      RECT 229.315 0.17 229.575 11.38 ;
      RECT 228.805 0.17 229.065 17.1 ;
      RECT 228.065 73.345 228.265 74.075 ;
      RECT 228.565 73.345 228.765 74.075 ;
      RECT 229.06 73.345 229.26 74.075 ;
      RECT 229.88 73.345 230.08 74.075 ;
      RECT 230.375 73.345 230.575 74.075 ;
      RECT 230.875 73.345 231.075 74.075 ;
      RECT 231.375 73.345 231.575 74.075 ;
      RECT 231.87 73.345 232.07 74.075 ;
      RECT 232.69 73.345 232.89 74.075 ;
      RECT 233.185 73.345 233.385 74.075 ;
      RECT 233.685 73.345 233.885 74.075 ;
      RECT 234.185 73.345 234.385 74.075 ;
      RECT 234.68 73.345 234.88 74.075 ;
      RECT 235.5 73.345 235.7 74.075 ;
      RECT 236.495 37.065 236.695 74.075 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 0 0.52 236.8 74.1 ;
      RECT 228.46 0 236.8 74.1 ;
      RECT 223.05 0 226.15 74.1 ;
      RECT 221.52 0 222.27 74.1 ;
      RECT 205.98 0 220.74 74.1 ;
      RECT 200.57 0 203.67 74.1 ;
      RECT 199.04 0 199.79 74.1 ;
      RECT 183.5 0 198.26 74.1 ;
      RECT 178.09 0 181.19 74.1 ;
      RECT 176.56 0 177.31 74.1 ;
      RECT 161.02 0 175.78 74.1 ;
      RECT 155.61 0 158.71 74.1 ;
      RECT 154.08 0 154.83 74.1 ;
      RECT 135 0.17 153.3 74.1 ;
      RECT 135.01 0 153.3 74.1 ;
      RECT 125.31 0 134.23 74.1 ;
      RECT 119.71 0 120.97 74.1 ;
      RECT 118.18 0 118.42 74.1 ;
      RECT 116.65 0 116.89 74.1 ;
      RECT 113.59 0 113.83 74.1 ;
      RECT 112.06 0 112.3 74.1 ;
      RECT 103.38 0 110.77 74.1 ;
      RECT 101.85 0 102.11 74.1 ;
      RECT 100.33 0 101.08 74.1 ;
      RECT 83.5 0 99.56 74.1 ;
      RECT 81.97 0 82.72 74.1 ;
      RECT 78.09 0 81.19 74.1 ;
      RECT 61.02 0 75.78 74.1 ;
      RECT 59.49 0 60.24 74.1 ;
      RECT 55.61 0 58.71 74.1 ;
      RECT 38.54 0 53.3 74.1 ;
      RECT 37.01 0 37.76 74.1 ;
      RECT 33.13 0 36.23 74.1 ;
      RECT 16.06 0 30.82 74.1 ;
      RECT 14.53 0 15.28 74.1 ;
      RECT 10.65 0 13.75 74.1 ;
      RECT 0 0 8.34 74.1 ;
    LAYER Metal3 ;
      RECT 0 0 236.8 74.1 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 138.09 0 145.17 74.1 ;
      RECT 132.94 0 134.76 74.1 ;
      RECT 127.79 0 129.61 74.1 ;
      RECT 232.8 0 236.8 74.1 ;
      RECT 227.18 0 229.47 74.1 ;
      RECT 227.18 30.685 236.8 36.805 ;
      RECT 221.56 0 223.85 74.1 ;
      RECT 215.94 0 218.23 74.1 ;
      RECT 215.94 30.685 223.85 36.805 ;
      RECT 210.32 0 212.61 74.1 ;
      RECT 204.7 0 206.99 74.1 ;
      RECT 204.7 30.685 212.61 36.805 ;
      RECT 199.08 0 201.37 74.1 ;
      RECT 193.46 0 195.75 74.1 ;
      RECT 193.46 30.685 201.37 36.805 ;
      RECT 187.84 0 190.13 74.1 ;
      RECT 52.29 0 54.58 74.1 ;
      RECT 46.67 0 48.96 74.1 ;
      RECT 46.67 30.685 54.58 36.805 ;
      RECT 41.05 0 43.34 74.1 ;
      RECT 35.43 0 37.72 74.1 ;
      RECT 35.43 30.685 43.34 36.805 ;
      RECT 29.81 0 32.1 74.1 ;
      RECT 24.19 0 26.48 74.1 ;
      RECT 24.19 30.685 32.1 36.805 ;
      RECT 18.57 0 20.86 74.1 ;
      RECT 12.95 0 15.24 74.1 ;
      RECT 12.95 30.685 20.86 36.805 ;
      RECT 7.33 0 9.62 74.1 ;
      RECT 0 0 4 74.1 ;
      RECT 0 30.685 9.62 36.805 ;
      RECT 182.22 0 184.51 74.1 ;
      RECT 182.22 30.685 190.13 36.805 ;
      RECT 176.6 0 178.89 74.1 ;
      RECT 170.98 0 173.27 74.1 ;
      RECT 170.98 30.685 178.89 36.805 ;
      RECT 165.36 0 167.65 74.1 ;
      RECT 159.74 0 162.03 74.1 ;
      RECT 159.74 30.685 167.65 36.805 ;
      RECT 154.12 0 156.41 74.1 ;
      RECT 148.5 0 150.79 74.1 ;
      RECT 148.5 30.685 156.41 36.805 ;
      RECT 122.64 0 124.46 74.1 ;
      RECT 117.49 0 119.31 74.1 ;
      RECT 112.34 0 114.16 74.1 ;
      RECT 107.19 0 109.01 74.1 ;
      RECT 102.04 0 103.86 74.1 ;
      RECT 91.63 0 98.71 74.1 ;
      RECT 86.01 0 88.3 74.1 ;
      RECT 80.39 0 82.68 74.1 ;
      RECT 80.39 30.685 88.3 36.805 ;
      RECT 74.77 0 77.06 74.1 ;
      RECT 69.15 0 71.44 74.1 ;
      RECT 69.15 30.685 77.06 36.805 ;
      RECT 63.53 0 65.82 74.1 ;
      RECT 57.91 0 60.2 74.1 ;
      RECT 57.91 30.685 65.82 36.805 ;
  END
END RM_IHPSG13_1P_256x8_c3_bm_bist

END LIBRARY
