# ------------------------------------------------------
#
#		Copyright 2025 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Wed Aug 27 13:14:43 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_256x32_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_256x32_c2_bm_bist 0 0 ;
  SIZE 702.83 BY 136.97 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 425.49 0 425.75 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.08 0 277.34 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 426 0 426.26 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.57 0 276.83 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 434.16 0 434.42 0.26 ;
    END
  END A_BM[16]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 268.41 0 268.67 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 432.785 0 433.045 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 269.785 0 270.045 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 418.35 0 418.61 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.22 0 284.48 0.26 ;
    END
  END A_DOUT[15]
  PIN B_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 428.04 0 428.3 0.26 ;
    END
  END B_DIN[16]
  PIN B_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 274.53 0 274.79 0.26 ;
    END
  END B_DIN[15]
  PIN B_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 426.51 0 426.77 0.26 ;
    END
  END B_BIST_DIN[16]
  PIN B_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 276.06 0 276.32 0.26 ;
    END
  END B_BIST_DIN[15]
  PIN B_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 419.525 0 419.785 0.26 ;
    END
  END B_BM[16]
  PIN B_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 283.045 0 283.305 0.26 ;
    END
  END B_BM[15]
  PIN B_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 421.055 0 421.315 0.26 ;
    END
  END B_BIST_BM[16]
  PIN B_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 281.515 0 281.775 0.26 ;
    END
  END B_BIST_BM[15]
  PIN B_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 435.18 0 435.44 0.26 ;
    END
  END B_DOUT[16]
  PIN B_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.39 0 267.65 0.26 ;
    END
  END B_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 683.425 0 687.845 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 665.745 0 670.165 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.065 0 652.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 630.385 0 634.805 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 612.705 0 617.125 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.025 0 599.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 577.345 0 581.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.665 0 564.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 541.985 0 546.405 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.305 0 528.725 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.625 0 511.045 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.945 0 493.365 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 471.265 0 475.685 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 453.585 0 458.005 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 435.905 0 440.325 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 418.225 0 422.645 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 388.635 0 391.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 378.335 0 381.145 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.885 0 365.695 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.585 0 355.395 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.435 0 350.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 337.135 0 339.945 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 321.685 0 324.495 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 311.385 0 314.195 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.185 0 284.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.505 0 266.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 244.825 0 249.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 227.145 0 231.565 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.465 0 213.885 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 191.785 0 196.205 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.105 0 178.525 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.425 0 160.845 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.745 0 143.165 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.065 0 125.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.385 0 107.805 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.705 0 90.125 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 136.97 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 692.265 0 696.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 674.585 0 679.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.905 0 661.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.225 0 643.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.545 0 625.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 603.865 0 608.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.185 0 590.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.505 0 572.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.825 0 555.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.145 0 537.565 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.465 0 519.885 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 497.785 0 502.205 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.105 0 484.525 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.425 0 466.845 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 444.745 0 449.165 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.065 0 431.485 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 383.485 0 386.295 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 373.185 0 375.995 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.035 0 370.845 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 357.735 0 360.545 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.285 0 345.095 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 331.985 0 334.795 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.835 0 329.645 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 316.535 0 319.345 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 0 275.765 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 0 258.085 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 0 240.405 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 0 222.725 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 0 205.045 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 0 187.365 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 0 169.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 0 152.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 0 134.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 0 116.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 0 98.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 0 81.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 692.265 53.41 696.685 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 674.585 53.41 679.005 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.905 53.41 661.325 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.225 53.41 643.645 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.545 53.41 625.965 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 603.865 53.41 608.285 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.185 53.41 590.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.505 53.41 572.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.825 53.41 555.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.145 53.41 537.565 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.465 53.41 519.885 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 497.785 53.41 502.205 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.105 53.41 484.525 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.425 53.41 466.845 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 444.745 53.41 449.165 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.065 53.41 431.485 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 53.41 275.765 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 53.41 258.085 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 53.41 240.405 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 53.41 222.725 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 53.41 205.045 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 53.41 187.365 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 53.41 169.685 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 53.41 152.005 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 53.41 134.325 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 53.41 116.645 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 53.41 98.965 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 53.41 81.285 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 136.97 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 136.97 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 443.17 0 443.43 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.4 0 259.66 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 443.68 0 443.94 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.89 0 259.15 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 451.84 0 452.1 0.26 ;
    END
  END A_BM[17]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 250.73 0 250.99 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 450.465 0 450.725 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 252.105 0 252.365 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 436.03 0 436.29 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.54 0 266.8 0.26 ;
    END
  END A_DOUT[14]
  PIN B_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 445.72 0 445.98 0.26 ;
    END
  END B_DIN[17]
  PIN B_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 256.85 0 257.11 0.26 ;
    END
  END B_DIN[14]
  PIN B_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 444.19 0 444.45 0.26 ;
    END
  END B_BIST_DIN[17]
  PIN B_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.38 0 258.64 0.26 ;
    END
  END B_BIST_DIN[14]
  PIN B_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 437.205 0 437.465 0.26 ;
    END
  END B_BM[17]
  PIN B_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 265.365 0 265.625 0.26 ;
    END
  END B_BM[14]
  PIN B_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 438.735 0 438.995 0.26 ;
    END
  END B_BIST_BM[17]
  PIN B_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 263.835 0 264.095 0.26 ;
    END
  END B_BIST_BM[14]
  PIN B_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 452.86 0 453.12 0.26 ;
    END
  END B_DOUT[17]
  PIN B_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.71 0 249.97 0.26 ;
    END
  END B_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 460.85 0 461.11 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.72 0 241.98 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.36 0 461.62 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.21 0 241.47 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 469.52 0 469.78 0.26 ;
    END
  END A_BM[18]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 233.05 0 233.31 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 468.145 0 468.405 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 234.425 0 234.685 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 453.71 0 453.97 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.86 0 249.12 0.26 ;
    END
  END A_DOUT[13]
  PIN B_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 463.4 0 463.66 0.26 ;
    END
  END B_DIN[18]
  PIN B_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 239.17 0 239.43 0.26 ;
    END
  END B_DIN[13]
  PIN B_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.87 0 462.13 0.26 ;
    END
  END B_BIST_DIN[18]
  PIN B_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 240.7 0 240.96 0.26 ;
    END
  END B_BIST_DIN[13]
  PIN B_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 454.885 0 455.145 0.26 ;
    END
  END B_BM[18]
  PIN B_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 247.685 0 247.945 0.26 ;
    END
  END B_BM[13]
  PIN B_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 456.415 0 456.675 0.26 ;
    END
  END B_BIST_BM[18]
  PIN B_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 246.155 0 246.415 0.26 ;
    END
  END B_BIST_BM[13]
  PIN B_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 470.54 0 470.8 0.26 ;
    END
  END B_DOUT[18]
  PIN B_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.03 0 232.29 0.26 ;
    END
  END B_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 478.53 0 478.79 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.04 0 224.3 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 479.04 0 479.3 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.53 0 223.79 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 487.2 0 487.46 0.26 ;
    END
  END A_BM[19]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.37 0 215.63 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 485.825 0 486.085 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 216.745 0 217.005 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 471.39 0 471.65 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.18 0 231.44 0.26 ;
    END
  END A_DOUT[12]
  PIN B_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 481.08 0 481.34 0.26 ;
    END
  END B_DIN[19]
  PIN B_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221.49 0 221.75 0.26 ;
    END
  END B_DIN[12]
  PIN B_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 479.55 0 479.81 0.26 ;
    END
  END B_BIST_DIN[19]
  PIN B_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.02 0 223.28 0.26 ;
    END
  END B_BIST_DIN[12]
  PIN B_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 472.565 0 472.825 0.26 ;
    END
  END B_BM[19]
  PIN B_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 230.005 0 230.265 0.26 ;
    END
  END B_BM[12]
  PIN B_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 474.095 0 474.355 0.26 ;
    END
  END B_BIST_BM[19]
  PIN B_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.475 0 228.735 0.26 ;
    END
  END B_BIST_BM[12]
  PIN B_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 488.22 0 488.48 0.26 ;
    END
  END B_DOUT[19]
  PIN B_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.35 0 214.61 0.26 ;
    END
  END B_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 496.21 0 496.47 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.36 0 206.62 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 496.72 0 496.98 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.85 0 206.11 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 504.88 0 505.14 0.26 ;
    END
  END A_BM[20]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 197.69 0 197.95 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 503.505 0 503.765 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 199.065 0 199.325 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 489.07 0 489.33 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.5 0 213.76 0.26 ;
    END
  END A_DOUT[11]
  PIN B_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 498.76 0 499.02 0.26 ;
    END
  END B_DIN[20]
  PIN B_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.81 0 204.07 0.26 ;
    END
  END B_DIN[11]
  PIN B_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 497.23 0 497.49 0.26 ;
    END
  END B_BIST_DIN[20]
  PIN B_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.34 0 205.6 0.26 ;
    END
  END B_BIST_DIN[11]
  PIN B_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 490.245 0 490.505 0.26 ;
    END
  END B_BM[20]
  PIN B_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 212.325 0 212.585 0.26 ;
    END
  END B_BM[11]
  PIN B_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 491.775 0 492.035 0.26 ;
    END
  END B_BIST_BM[20]
  PIN B_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 210.795 0 211.055 0.26 ;
    END
  END B_BIST_BM[11]
  PIN B_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 505.9 0 506.16 0.26 ;
    END
  END B_DOUT[20]
  PIN B_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.67 0 196.93 0.26 ;
    END
  END B_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 513.89 0 514.15 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.68 0 188.94 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.4 0 514.66 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.17 0 188.43 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 522.56 0 522.82 0.26 ;
    END
  END A_BM[21]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 180.01 0 180.27 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 521.185 0 521.445 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 181.385 0 181.645 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 506.75 0 507.01 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.82 0 196.08 0.26 ;
    END
  END A_DOUT[10]
  PIN B_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 516.44 0 516.7 0.26 ;
    END
  END B_DIN[21]
  PIN B_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 186.13 0 186.39 0.26 ;
    END
  END B_DIN[10]
  PIN B_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.91 0 515.17 0.26 ;
    END
  END B_BIST_DIN[21]
  PIN B_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 187.66 0 187.92 0.26 ;
    END
  END B_BIST_DIN[10]
  PIN B_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 507.925 0 508.185 0.26 ;
    END
  END B_BM[21]
  PIN B_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 194.645 0 194.905 0.26 ;
    END
  END B_BM[10]
  PIN B_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 509.455 0 509.715 0.26 ;
    END
  END B_BIST_BM[21]
  PIN B_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.115 0 193.375 0.26 ;
    END
  END B_BIST_BM[10]
  PIN B_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 523.58 0 523.84 0.26 ;
    END
  END B_DOUT[21]
  PIN B_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.99 0 179.25 0.26 ;
    END
  END B_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 531.57 0 531.83 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171 0 171.26 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 532.08 0 532.34 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 170.49 0 170.75 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 540.24 0 540.5 0.26 ;
    END
  END A_BM[22]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 162.33 0 162.59 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 538.865 0 539.125 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 163.705 0 163.965 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 524.43 0 524.69 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.14 0 178.4 0.26 ;
    END
  END A_DOUT[9]
  PIN B_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 534.12 0 534.38 0.26 ;
    END
  END B_DIN[22]
  PIN B_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.45 0 168.71 0.26 ;
    END
  END B_DIN[9]
  PIN B_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 532.59 0 532.85 0.26 ;
    END
  END B_BIST_DIN[22]
  PIN B_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 169.98 0 170.24 0.26 ;
    END
  END B_BIST_DIN[9]
  PIN B_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 525.605 0 525.865 0.26 ;
    END
  END B_BM[22]
  PIN B_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.965 0 177.225 0.26 ;
    END
  END B_BM[9]
  PIN B_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 527.135 0 527.395 0.26 ;
    END
  END B_BIST_BM[22]
  PIN B_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 175.435 0 175.695 0.26 ;
    END
  END B_BIST_BM[9]
  PIN B_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 541.26 0 541.52 0.26 ;
    END
  END B_DOUT[22]
  PIN B_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.31 0 161.57 0.26 ;
    END
  END B_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 549.25 0 549.51 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.32 0 153.58 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 549.76 0 550.02 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.81 0 153.07 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 557.92 0 558.18 0.26 ;
    END
  END A_BM[23]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.65 0 144.91 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 556.545 0 556.805 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.025 0 146.285 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 542.11 0 542.37 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.46 0 160.72 0.26 ;
    END
  END A_DOUT[8]
  PIN B_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 551.8 0 552.06 0.26 ;
    END
  END B_DIN[23]
  PIN B_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.77 0 151.03 0.26 ;
    END
  END B_DIN[8]
  PIN B_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 550.27 0 550.53 0.26 ;
    END
  END B_BIST_DIN[23]
  PIN B_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 152.3 0 152.56 0.26 ;
    END
  END B_BIST_DIN[8]
  PIN B_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 543.285 0 543.545 0.26 ;
    END
  END B_BM[23]
  PIN B_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 159.285 0 159.545 0.26 ;
    END
  END B_BM[8]
  PIN B_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 544.815 0 545.075 0.26 ;
    END
  END B_BIST_BM[23]
  PIN B_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.755 0 158.015 0.26 ;
    END
  END B_BIST_BM[8]
  PIN B_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 558.94 0 559.2 0.26 ;
    END
  END B_DOUT[23]
  PIN B_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.63 0 143.89 0.26 ;
    END
  END B_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 566.93 0 567.19 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.64 0 135.9 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 567.44 0 567.7 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.13 0 135.39 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 575.6 0 575.86 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.97 0 127.23 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 574.225 0 574.485 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 128.345 0 128.605 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 559.79 0 560.05 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.78 0 143.04 0.26 ;
    END
  END A_DOUT[7]
  PIN B_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 569.48 0 569.74 0.26 ;
    END
  END B_DIN[24]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.09 0 133.35 0.26 ;
    END
  END B_DIN[7]
  PIN B_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 567.95 0 568.21 0.26 ;
    END
  END B_BIST_DIN[24]
  PIN B_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.62 0 134.88 0.26 ;
    END
  END B_BIST_DIN[7]
  PIN B_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 560.965 0 561.225 0.26 ;
    END
  END B_BM[24]
  PIN B_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 141.605 0 141.865 0.26 ;
    END
  END B_BM[7]
  PIN B_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 562.495 0 562.755 0.26 ;
    END
  END B_BIST_BM[24]
  PIN B_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 140.075 0 140.335 0.26 ;
    END
  END B_BIST_BM[7]
  PIN B_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 576.62 0 576.88 0.26 ;
    END
  END B_DOUT[24]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.95 0 126.21 0.26 ;
    END
  END B_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 584.61 0 584.87 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.96 0 118.22 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.12 0 585.38 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.45 0 117.71 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 593.28 0 593.54 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.29 0 109.55 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 591.905 0 592.165 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.665 0 110.925 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 577.47 0 577.73 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.1 0 125.36 0.26 ;
    END
  END A_DOUT[6]
  PIN B_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 587.16 0 587.42 0.26 ;
    END
  END B_DIN[25]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.41 0 115.67 0.26 ;
    END
  END B_DIN[6]
  PIN B_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.63 0 585.89 0.26 ;
    END
  END B_BIST_DIN[25]
  PIN B_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.94 0 117.2 0.26 ;
    END
  END B_BIST_DIN[6]
  PIN B_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 578.645 0 578.905 0.26 ;
    END
  END B_BM[25]
  PIN B_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.925 0 124.185 0.26 ;
    END
  END B_BM[6]
  PIN B_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 580.175 0 580.435 0.26 ;
    END
  END B_BIST_BM[25]
  PIN B_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.395 0 122.655 0.26 ;
    END
  END B_BIST_BM[6]
  PIN B_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 594.3 0 594.56 0.26 ;
    END
  END B_DOUT[25]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.27 0 108.53 0.26 ;
    END
  END B_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 602.29 0 602.55 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.28 0 100.54 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 602.8 0 603.06 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.77 0 100.03 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 610.96 0 611.22 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 91.61 0 91.87 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 609.585 0 609.845 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 92.985 0 93.245 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 595.15 0 595.41 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 107.42 0 107.68 0.26 ;
    END
  END A_DOUT[5]
  PIN B_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 604.84 0 605.1 0.26 ;
    END
  END B_DIN[26]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 97.73 0 97.99 0.26 ;
    END
  END B_DIN[5]
  PIN B_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 603.31 0 603.57 0.26 ;
    END
  END B_BIST_DIN[26]
  PIN B_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.26 0 99.52 0.26 ;
    END
  END B_BIST_DIN[5]
  PIN B_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 596.325 0 596.585 0.26 ;
    END
  END B_BM[26]
  PIN B_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 106.245 0 106.505 0.26 ;
    END
  END B_BM[5]
  PIN B_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 597.855 0 598.115 0.26 ;
    END
  END B_BIST_BM[26]
  PIN B_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.715 0 104.975 0.26 ;
    END
  END B_BIST_BM[5]
  PIN B_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 611.98 0 612.24 0.26 ;
    END
  END B_DOUT[26]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 90.59 0 90.85 0.26 ;
    END
  END B_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 619.97 0 620.23 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.6 0 82.86 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 620.48 0 620.74 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.09 0 82.35 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 628.64 0 628.9 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 73.93 0 74.19 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 627.265 0 627.525 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 75.305 0 75.565 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 612.83 0 613.09 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.74 0 90 0.26 ;
    END
  END A_DOUT[4]
  PIN B_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 622.52 0 622.78 0.26 ;
    END
  END B_DIN[27]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 80.05 0 80.31 0.26 ;
    END
  END B_DIN[4]
  PIN B_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 620.99 0 621.25 0.26 ;
    END
  END B_BIST_DIN[27]
  PIN B_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.58 0 81.84 0.26 ;
    END
  END B_BIST_DIN[4]
  PIN B_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 614.005 0 614.265 0.26 ;
    END
  END B_BM[27]
  PIN B_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.565 0 88.825 0.26 ;
    END
  END B_BM[4]
  PIN B_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 615.535 0 615.795 0.26 ;
    END
  END B_BIST_BM[27]
  PIN B_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 87.035 0 87.295 0.26 ;
    END
  END B_BIST_BM[4]
  PIN B_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 629.66 0 629.92 0.26 ;
    END
  END B_DOUT[27]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.91 0 73.17 0.26 ;
    END
  END B_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 637.65 0 637.91 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 638.16 0 638.42 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.41 0 64.67 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 646.32 0 646.58 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.25 0 56.51 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 644.945 0 645.205 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.625 0 57.885 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 630.51 0 630.77 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 640.2 0 640.46 0.26 ;
    END
  END B_DIN[28]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 638.67 0 638.93 0.26 ;
    END
  END B_BIST_DIN[28]
  PIN B_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 63.9 0 64.16 0.26 ;
    END
  END B_BIST_DIN[3]
  PIN B_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 631.685 0 631.945 0.26 ;
    END
  END B_BM[28]
  PIN B_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.885 0 71.145 0.26 ;
    END
  END B_BM[3]
  PIN B_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 633.215 0 633.475 0.26 ;
    END
  END B_BIST_BM[28]
  PIN B_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.355 0 69.615 0.26 ;
    END
  END B_BIST_BM[3]
  PIN B_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 647.34 0 647.6 0.26 ;
    END
  END B_DOUT[28]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 655.33 0 655.59 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 655.84 0 656.1 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.73 0 46.99 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 664 0 664.26 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.57 0 38.83 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 662.625 0 662.885 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 39.945 0 40.205 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 648.19 0 648.45 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 657.88 0 658.14 0.26 ;
    END
  END B_DIN[29]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 656.35 0 656.61 0.26 ;
    END
  END B_BIST_DIN[29]
  PIN B_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 46.22 0 46.48 0.26 ;
    END
  END B_BIST_DIN[2]
  PIN B_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 649.365 0 649.625 0.26 ;
    END
  END B_BM[29]
  PIN B_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.205 0 53.465 0.26 ;
    END
  END B_BM[2]
  PIN B_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 650.895 0 651.155 0.26 ;
    END
  END B_BIST_BM[29]
  PIN B_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 51.675 0 51.935 0.26 ;
    END
  END B_BIST_BM[2]
  PIN B_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 665.02 0 665.28 0.26 ;
    END
  END B_DOUT[29]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 673.01 0 673.27 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 673.52 0 673.78 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.05 0 29.31 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 681.68 0 681.94 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.89 0 21.15 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 680.305 0 680.565 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.265 0 22.525 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 665.87 0 666.13 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 675.56 0 675.82 0.26 ;
    END
  END B_DIN[30]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 674.03 0 674.29 0.26 ;
    END
  END B_BIST_DIN[30]
  PIN B_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 28.54 0 28.8 0.26 ;
    END
  END B_BIST_DIN[1]
  PIN B_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 667.045 0 667.305 0.26 ;
    END
  END B_BM[30]
  PIN B_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 35.525 0 35.785 0.26 ;
    END
  END B_BM[1]
  PIN B_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 668.575 0 668.835 0.26 ;
    END
  END B_BIST_BM[30]
  PIN B_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.995 0 34.255 0.26 ;
    END
  END B_BIST_BM[1]
  PIN B_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 682.7 0 682.96 0.26 ;
    END
  END B_DOUT[30]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 690.69 0 690.95 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 691.2 0 691.46 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.136375 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.874907 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.37 0 11.63 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 699.36 0 699.62 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7264 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.501618 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.21 0 3.47 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 697.985 0 698.245 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7602 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.678367 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.585 0 4.845 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 683.55 0 683.81 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 693.24 0 693.5 0.26 ;
    END
  END B_DIN[31]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 691.71 0 691.97 0.26 ;
    END
  END B_BIST_DIN[31]
  PIN B_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9445 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.929052 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.86 0 11.12 0.26 ;
    END
  END B_BIST_DIN[0]
  PIN B_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 684.725 0 684.985 0.26 ;
    END
  END B_BM[31]
  PIN B_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 17.845 0 18.105 0.26 ;
    END
  END B_BM[0]
  PIN B_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 686.255 0 686.515 0.26 ;
    END
  END B_BIST_BM[31]
  PIN B_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 16.315 0 16.575 0.26 ;
    END
  END B_BIST_BM[0]
  PIN B_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 700.38 0 700.64 0.26 ;
    END
  END B_DOUT[31]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 367.505 0 367.765 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.115 0 373.375 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 335.065 0 335.325 0.26 ;
    END
  END B_ADDR[0]
  PIN B_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8293 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.84466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 329.455 0 329.715 0.26 ;
    END
  END B_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.015 0 368.275 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 373.625 0 373.885 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.555 0 334.815 0.26 ;
    END
  END B_ADDR[1]
  PIN B_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1459 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.378641 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 328.945 0 329.205 0.26 ;
    END
  END B_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 376.685 0 376.945 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 377.195 0 377.455 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 325.885 0 326.145 0.26 ;
    END
  END B_ADDR[2]
  PIN B_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 325.375 0 325.635 0.26 ;
    END
  END B_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 375.665 0 375.925 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 376.175 0 376.435 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 326.905 0 327.165 0.26 ;
    END
  END B_ADDR[3]
  PIN B_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.7317 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.935524 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 326.395 0 326.655 0.26 ;
    END
  END B_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.285 0 356.545 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.795 0 357.055 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.285 0 346.545 0.26 ;
    END
  END B_ADDR[4]
  PIN B_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4677 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.938511 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 345.775 0 346.035 0.26 ;
    END
  END B_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.265 0 355.525 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.775 0 356.035 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.305 0 347.565 0.26 ;
    END
  END B_ADDR[5]
  PIN B_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9937 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 65.599701 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.795 0 347.055 0.26 ;
    END
  END B_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.235 0 379.495 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.725 0 378.985 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN B_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3819 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 72.511327 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 323.335 0 323.595 0.26 ;
    END
  END B_ADDR[6]
  PIN B_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1167 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 71.190939 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 323.845 0 324.105 0.26 ;
    END
  END B_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.215 0 378.475 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 377.705 0 377.965 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN B_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3761 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 82.440129 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 324.355 0 324.615 0.26 ;
    END
  END B_ADDR[7]
  PIN B_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1109 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 81.119741 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 324.865 0 325.125 0.26 ;
    END
  END B_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 365.975 0 366.235 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.545 0 369.805 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.035 0 369.295 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 366.485 0 366.745 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 386.885 0 387.145 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 336.595 0 336.855 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.025 0 333.285 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.535 0 333.795 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 336.085 0 336.345 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.685 0 315.945 0.26 ;
    END
  END B_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 258.2003 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.17 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.266993 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.674515 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.525 0 368.785 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.445 0 364.705 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.075 0 371.335 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 370.565 0 370.825 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.955 0 365.215 0.26 ;
    END
  END A_BIST_MEN
  PIN B_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 258.7774 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 27.17 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.197902 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.695755 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.045 0 334.305 0.26 ;
    END
  END B_BIST_EN
  PIN B_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.125 0 338.385 0.26 ;
    END
  END B_BIST_CLK
  PIN B_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 331.495 0 331.755 0.26 ;
    END
  END B_BIST_REN
  PIN B_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 332.005 0 332.265 0.26 ;
    END
  END B_BIST_WEN
  PIN B_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.615 0 337.875 0.26 ;
    END
  END B_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 702.83 136.97 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 136.94 ;
      RECT 1.135 136.21 1.335 136.94 ;
      RECT 1.545 136.21 1.905 136.94 ;
      RECT 2.115 136.21 2.315 136.94 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 136.21 2.97 136.94 ;
      RECT 3.21 0.52 3.47 5.57 ;
      RECT 3.18 136.21 3.54 136.94 ;
      RECT 3.835 136.21 4.035 136.94 ;
      RECT 4.33 136.21 4.69 136.94 ;
      RECT 4.585 0.52 4.845 6.28 ;
      RECT 4.9 136.21 5.1 136.94 ;
      RECT 5.555 136.21 5.755 136.94 ;
      RECT 5.965 136.21 6.325 136.94 ;
      RECT 6.535 136.21 6.735 136.94 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 136.21 7.39 136.94 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 136.21 7.96 136.94 ;
      RECT 8.255 136.21 8.455 136.94 ;
      RECT 8.75 136.21 9.11 136.94 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 136.21 9.52 136.94 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 136.21 10.175 136.94 ;
      RECT 10.385 136.21 10.745 136.94 ;
      RECT 10.86 0.52 11.12 11.315 ;
      RECT 10.955 136.21 11.155 136.94 ;
      RECT 11.37 0.52 11.63 13.45 ;
      RECT 11.61 136.21 11.81 136.94 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 136.21 12.38 136.94 ;
      RECT 12.675 136.21 12.875 136.94 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 136.21 13.53 136.94 ;
      RECT 13.74 136.21 13.94 136.94 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 136.21 14.595 136.94 ;
      RECT 14.805 136.21 15.165 136.94 ;
      RECT 15.375 136.21 15.575 136.94 ;
      RECT 16.03 136.21 16.23 136.94 ;
      RECT 16.315 0.52 16.575 2.82 ;
      RECT 16.44 136.21 16.8 136.94 ;
      RECT 17.095 136.21 17.295 136.94 ;
      RECT 17.59 136.21 17.95 136.94 ;
      RECT 17.845 0.52 18.105 2.82 ;
      RECT 18.16 136.21 18.36 136.94 ;
      RECT 18.815 136.21 19.015 136.94 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 136.21 19.585 136.94 ;
      RECT 19.795 136.21 19.995 136.94 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 136.21 20.65 136.94 ;
      RECT 20.89 0.52 21.15 5.57 ;
      RECT 20.86 136.21 21.22 136.94 ;
      RECT 21.515 136.21 21.715 136.94 ;
      RECT 22.01 136.21 22.37 136.94 ;
      RECT 22.265 0.52 22.525 6.28 ;
      RECT 22.58 136.21 22.78 136.94 ;
      RECT 23.235 136.21 23.435 136.94 ;
      RECT 23.645 136.21 24.005 136.94 ;
      RECT 24.215 136.21 24.415 136.94 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 136.21 25.07 136.94 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 136.21 25.64 136.94 ;
      RECT 25.935 136.21 26.135 136.94 ;
      RECT 26.43 136.21 26.79 136.94 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 136.21 27.2 136.94 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 136.21 27.855 136.94 ;
      RECT 28.065 136.21 28.425 136.94 ;
      RECT 28.54 0.52 28.8 11.315 ;
      RECT 28.635 136.21 28.835 136.94 ;
      RECT 29.05 0.52 29.31 13.45 ;
      RECT 29.29 136.21 29.49 136.94 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 136.21 30.06 136.94 ;
      RECT 30.355 136.21 30.555 136.94 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 136.21 31.21 136.94 ;
      RECT 31.42 136.21 31.62 136.94 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 136.21 32.275 136.94 ;
      RECT 32.485 136.21 32.845 136.94 ;
      RECT 33.055 136.21 33.255 136.94 ;
      RECT 33.71 136.21 33.91 136.94 ;
      RECT 33.995 0.52 34.255 2.82 ;
      RECT 34.12 136.21 34.48 136.94 ;
      RECT 34.775 136.21 34.975 136.94 ;
      RECT 35.27 136.21 35.63 136.94 ;
      RECT 35.525 0.52 35.785 2.82 ;
      RECT 35.84 136.21 36.04 136.94 ;
      RECT 36.495 136.21 36.695 136.94 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 136.21 37.265 136.94 ;
      RECT 37.475 136.21 37.675 136.94 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 136.21 38.33 136.94 ;
      RECT 38.57 0.52 38.83 5.57 ;
      RECT 38.54 136.21 38.9 136.94 ;
      RECT 39.195 136.21 39.395 136.94 ;
      RECT 39.69 136.21 40.05 136.94 ;
      RECT 39.945 0.52 40.205 6.28 ;
      RECT 40.26 136.21 40.46 136.94 ;
      RECT 40.915 136.21 41.115 136.94 ;
      RECT 41.325 136.21 41.685 136.94 ;
      RECT 41.895 136.21 42.095 136.94 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 136.21 42.75 136.94 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 136.21 43.32 136.94 ;
      RECT 43.615 136.21 43.815 136.94 ;
      RECT 44.11 136.21 44.47 136.94 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 136.21 44.88 136.94 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 136.21 45.535 136.94 ;
      RECT 45.745 136.21 46.105 136.94 ;
      RECT 46.22 0.52 46.48 11.315 ;
      RECT 46.315 136.21 46.515 136.94 ;
      RECT 46.73 0.52 46.99 13.45 ;
      RECT 46.97 136.21 47.17 136.94 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 136.21 47.74 136.94 ;
      RECT 48.035 136.21 48.235 136.94 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 136.21 48.89 136.94 ;
      RECT 49.1 136.21 49.3 136.94 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 136.21 49.955 136.94 ;
      RECT 50.165 136.21 50.525 136.94 ;
      RECT 50.735 136.21 50.935 136.94 ;
      RECT 51.39 136.21 51.59 136.94 ;
      RECT 51.675 0.52 51.935 2.82 ;
      RECT 51.8 136.21 52.16 136.94 ;
      RECT 52.455 136.21 52.655 136.94 ;
      RECT 52.95 136.21 53.31 136.94 ;
      RECT 53.205 0.52 53.465 2.82 ;
      RECT 53.52 136.21 53.72 136.94 ;
      RECT 54.175 136.21 54.375 136.94 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 136.21 54.945 136.94 ;
      RECT 55.155 136.21 55.355 136.94 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 136.21 56.01 136.94 ;
      RECT 56.25 0.52 56.51 5.57 ;
      RECT 56.22 136.21 56.58 136.94 ;
      RECT 56.875 136.21 57.075 136.94 ;
      RECT 57.37 136.21 57.73 136.94 ;
      RECT 57.625 0.52 57.885 6.28 ;
      RECT 57.94 136.21 58.14 136.94 ;
      RECT 58.595 136.21 58.795 136.94 ;
      RECT 59.005 136.21 59.365 136.94 ;
      RECT 59.575 136.21 59.775 136.94 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 136.21 60.43 136.94 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 136.21 61 136.94 ;
      RECT 61.295 136.21 61.495 136.94 ;
      RECT 61.79 136.21 62.15 136.94 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 136.21 62.56 136.94 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 136.21 63.215 136.94 ;
      RECT 63.425 136.21 63.785 136.94 ;
      RECT 63.9 0.52 64.16 11.315 ;
      RECT 63.995 136.21 64.195 136.94 ;
      RECT 64.41 0.52 64.67 13.45 ;
      RECT 64.65 136.21 64.85 136.94 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 136.21 65.42 136.94 ;
      RECT 65.715 136.21 65.915 136.94 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 136.21 66.57 136.94 ;
      RECT 66.78 136.21 66.98 136.94 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 136.21 67.635 136.94 ;
      RECT 67.845 136.21 68.205 136.94 ;
      RECT 68.415 136.21 68.615 136.94 ;
      RECT 69.07 136.21 69.27 136.94 ;
      RECT 69.355 0.52 69.615 2.82 ;
      RECT 69.48 136.21 69.84 136.94 ;
      RECT 70.135 136.21 70.335 136.94 ;
      RECT 70.63 136.21 70.99 136.94 ;
      RECT 70.885 0.52 71.145 2.82 ;
      RECT 71.2 136.21 71.4 136.94 ;
      RECT 71.855 136.21 72.055 136.94 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 72.265 136.21 72.625 136.94 ;
      RECT 72.835 136.21 73.035 136.94 ;
      RECT 72.91 0.52 73.17 7.78 ;
      RECT 73.42 0.3 73.68 5.235 ;
      RECT 73.49 136.21 73.69 136.94 ;
      RECT 73.93 0.52 74.19 5.57 ;
      RECT 73.9 136.21 74.26 136.94 ;
      RECT 74.555 136.21 74.755 136.94 ;
      RECT 75.05 136.21 75.41 136.94 ;
      RECT 75.305 0.52 75.565 6.28 ;
      RECT 75.62 136.21 75.82 136.94 ;
      RECT 76.275 136.21 76.475 136.94 ;
      RECT 76.685 136.21 77.045 136.94 ;
      RECT 77.255 136.21 77.455 136.94 ;
      RECT 76.99 0.18 77.76 0.88 ;
      RECT 77.91 136.21 78.11 136.94 ;
      RECT 78.01 0.3 78.27 8.7 ;
      RECT 78.32 136.21 78.68 136.94 ;
      RECT 78.975 136.21 79.175 136.94 ;
      RECT 79.47 136.21 79.83 136.94 ;
      RECT 80.56 0.155 81.33 0.445 ;
      RECT 80.56 0.155 80.82 8.665 ;
      RECT 81.07 0.155 81.33 8.665 ;
      RECT 80.04 136.21 80.24 136.94 ;
      RECT 80.05 0.52 80.31 9.955 ;
      RECT 80.695 136.21 80.895 136.94 ;
      RECT 81.105 136.21 81.465 136.94 ;
      RECT 81.58 0.52 81.84 11.315 ;
      RECT 81.675 136.21 81.875 136.94 ;
      RECT 82.09 0.52 82.35 13.45 ;
      RECT 82.33 136.21 82.53 136.94 ;
      RECT 82.6 0.52 82.86 14.115 ;
      RECT 82.74 136.21 83.1 136.94 ;
      RECT 83.395 136.21 83.595 136.94 ;
      RECT 84.795 0.155 85.565 0.445 ;
      RECT 84.795 0.155 85.055 13.21 ;
      RECT 85.305 0.155 85.565 13.21 ;
      RECT 83.89 136.21 84.25 136.94 ;
      RECT 84.46 136.21 84.66 136.94 ;
      RECT 85.815 0.18 86.585 0.88 ;
      RECT 85.815 0.18 86.075 12.9 ;
      RECT 86.325 0.18 86.585 12.9 ;
      RECT 85.115 136.21 85.315 136.94 ;
      RECT 85.525 136.21 85.885 136.94 ;
      RECT 86.095 136.21 86.295 136.94 ;
      RECT 86.75 136.21 86.95 136.94 ;
      RECT 87.035 0.52 87.295 2.82 ;
      RECT 87.16 136.21 87.52 136.94 ;
      RECT 87.815 136.21 88.015 136.94 ;
      RECT 88.31 136.21 88.67 136.94 ;
      RECT 88.565 0.52 88.825 2.82 ;
      RECT 88.88 136.21 89.08 136.94 ;
      RECT 89.535 136.21 89.735 136.94 ;
      RECT 89.74 0.52 90 4.315 ;
      RECT 89.945 136.21 90.305 136.94 ;
      RECT 90.515 136.21 90.715 136.94 ;
      RECT 90.59 0.52 90.85 7.78 ;
      RECT 91.1 0.3 91.36 5.235 ;
      RECT 91.17 136.21 91.37 136.94 ;
      RECT 91.61 0.52 91.87 5.57 ;
      RECT 91.58 136.21 91.94 136.94 ;
      RECT 92.235 136.21 92.435 136.94 ;
      RECT 92.73 136.21 93.09 136.94 ;
      RECT 92.985 0.52 93.245 6.28 ;
      RECT 93.3 136.21 93.5 136.94 ;
      RECT 93.955 136.21 94.155 136.94 ;
      RECT 94.365 136.21 94.725 136.94 ;
      RECT 94.935 136.21 95.135 136.94 ;
      RECT 94.67 0.18 95.44 0.88 ;
      RECT 95.59 136.21 95.79 136.94 ;
      RECT 95.69 0.3 95.95 8.7 ;
      RECT 96 136.21 96.36 136.94 ;
      RECT 96.655 136.21 96.855 136.94 ;
      RECT 97.15 136.21 97.51 136.94 ;
      RECT 98.24 0.155 99.01 0.445 ;
      RECT 98.24 0.155 98.5 8.665 ;
      RECT 98.75 0.155 99.01 8.665 ;
      RECT 97.72 136.21 97.92 136.94 ;
      RECT 97.73 0.52 97.99 9.955 ;
      RECT 98.375 136.21 98.575 136.94 ;
      RECT 98.785 136.21 99.145 136.94 ;
      RECT 99.26 0.52 99.52 11.315 ;
      RECT 99.355 136.21 99.555 136.94 ;
      RECT 99.77 0.52 100.03 13.45 ;
      RECT 100.01 136.21 100.21 136.94 ;
      RECT 100.28 0.52 100.54 14.115 ;
      RECT 100.42 136.21 100.78 136.94 ;
      RECT 101.075 136.21 101.275 136.94 ;
      RECT 102.475 0.155 103.245 0.445 ;
      RECT 102.475 0.155 102.735 13.21 ;
      RECT 102.985 0.155 103.245 13.21 ;
      RECT 101.57 136.21 101.93 136.94 ;
      RECT 102.14 136.21 102.34 136.94 ;
      RECT 103.495 0.18 104.265 0.88 ;
      RECT 103.495 0.18 103.755 12.9 ;
      RECT 104.005 0.18 104.265 12.9 ;
      RECT 102.795 136.21 102.995 136.94 ;
      RECT 103.205 136.21 103.565 136.94 ;
      RECT 103.775 136.21 103.975 136.94 ;
      RECT 104.43 136.21 104.63 136.94 ;
      RECT 104.715 0.52 104.975 2.82 ;
      RECT 104.84 136.21 105.2 136.94 ;
      RECT 105.495 136.21 105.695 136.94 ;
      RECT 105.99 136.21 106.35 136.94 ;
      RECT 106.245 0.52 106.505 2.82 ;
      RECT 106.56 136.21 106.76 136.94 ;
      RECT 107.215 136.21 107.415 136.94 ;
      RECT 107.42 0.52 107.68 4.315 ;
      RECT 107.625 136.21 107.985 136.94 ;
      RECT 108.195 136.21 108.395 136.94 ;
      RECT 108.27 0.52 108.53 7.78 ;
      RECT 108.78 0.3 109.04 5.235 ;
      RECT 108.85 136.21 109.05 136.94 ;
      RECT 109.29 0.52 109.55 5.57 ;
      RECT 109.26 136.21 109.62 136.94 ;
      RECT 109.915 136.21 110.115 136.94 ;
      RECT 110.41 136.21 110.77 136.94 ;
      RECT 110.665 0.52 110.925 6.28 ;
      RECT 110.98 136.21 111.18 136.94 ;
      RECT 111.635 136.21 111.835 136.94 ;
      RECT 112.045 136.21 112.405 136.94 ;
      RECT 112.615 136.21 112.815 136.94 ;
      RECT 112.35 0.18 113.12 0.88 ;
      RECT 113.27 136.21 113.47 136.94 ;
      RECT 113.37 0.3 113.63 8.7 ;
      RECT 113.68 136.21 114.04 136.94 ;
      RECT 114.335 136.21 114.535 136.94 ;
      RECT 114.83 136.21 115.19 136.94 ;
      RECT 115.92 0.155 116.69 0.445 ;
      RECT 115.92 0.155 116.18 8.665 ;
      RECT 116.43 0.155 116.69 8.665 ;
      RECT 115.4 136.21 115.6 136.94 ;
      RECT 115.41 0.52 115.67 9.955 ;
      RECT 116.055 136.21 116.255 136.94 ;
      RECT 116.465 136.21 116.825 136.94 ;
      RECT 116.94 0.52 117.2 11.315 ;
      RECT 117.035 136.21 117.235 136.94 ;
      RECT 117.45 0.52 117.71 13.45 ;
      RECT 117.69 136.21 117.89 136.94 ;
      RECT 117.96 0.52 118.22 14.115 ;
      RECT 118.1 136.21 118.46 136.94 ;
      RECT 118.755 136.21 118.955 136.94 ;
      RECT 120.155 0.155 120.925 0.445 ;
      RECT 120.155 0.155 120.415 13.21 ;
      RECT 120.665 0.155 120.925 13.21 ;
      RECT 119.25 136.21 119.61 136.94 ;
      RECT 119.82 136.21 120.02 136.94 ;
      RECT 121.175 0.18 121.945 0.88 ;
      RECT 121.175 0.18 121.435 12.9 ;
      RECT 121.685 0.18 121.945 12.9 ;
      RECT 120.475 136.21 120.675 136.94 ;
      RECT 120.885 136.21 121.245 136.94 ;
      RECT 121.455 136.21 121.655 136.94 ;
      RECT 122.11 136.21 122.31 136.94 ;
      RECT 122.395 0.52 122.655 2.82 ;
      RECT 122.52 136.21 122.88 136.94 ;
      RECT 123.175 136.21 123.375 136.94 ;
      RECT 123.67 136.21 124.03 136.94 ;
      RECT 123.925 0.52 124.185 2.82 ;
      RECT 124.24 136.21 124.44 136.94 ;
      RECT 124.895 136.21 125.095 136.94 ;
      RECT 125.1 0.52 125.36 4.315 ;
      RECT 125.305 136.21 125.665 136.94 ;
      RECT 125.875 136.21 126.075 136.94 ;
      RECT 125.95 0.52 126.21 7.78 ;
      RECT 126.46 0.3 126.72 5.235 ;
      RECT 126.53 136.21 126.73 136.94 ;
      RECT 126.97 0.52 127.23 5.57 ;
      RECT 126.94 136.21 127.3 136.94 ;
      RECT 127.595 136.21 127.795 136.94 ;
      RECT 128.09 136.21 128.45 136.94 ;
      RECT 128.345 0.52 128.605 6.28 ;
      RECT 128.66 136.21 128.86 136.94 ;
      RECT 129.315 136.21 129.515 136.94 ;
      RECT 129.725 136.21 130.085 136.94 ;
      RECT 130.295 136.21 130.495 136.94 ;
      RECT 130.03 0.18 130.8 0.88 ;
      RECT 130.95 136.21 131.15 136.94 ;
      RECT 131.05 0.3 131.31 8.7 ;
      RECT 131.36 136.21 131.72 136.94 ;
      RECT 132.015 136.21 132.215 136.94 ;
      RECT 132.51 136.21 132.87 136.94 ;
      RECT 133.6 0.155 134.37 0.445 ;
      RECT 133.6 0.155 133.86 8.665 ;
      RECT 134.11 0.155 134.37 8.665 ;
      RECT 133.08 136.21 133.28 136.94 ;
      RECT 133.09 0.52 133.35 9.955 ;
      RECT 133.735 136.21 133.935 136.94 ;
      RECT 134.145 136.21 134.505 136.94 ;
      RECT 134.62 0.52 134.88 11.315 ;
      RECT 134.715 136.21 134.915 136.94 ;
      RECT 135.13 0.52 135.39 13.45 ;
      RECT 135.37 136.21 135.57 136.94 ;
      RECT 135.64 0.52 135.9 14.115 ;
      RECT 135.78 136.21 136.14 136.94 ;
      RECT 136.435 136.21 136.635 136.94 ;
      RECT 137.835 0.155 138.605 0.445 ;
      RECT 137.835 0.155 138.095 13.21 ;
      RECT 138.345 0.155 138.605 13.21 ;
      RECT 136.93 136.21 137.29 136.94 ;
      RECT 137.5 136.21 137.7 136.94 ;
      RECT 138.855 0.18 139.625 0.88 ;
      RECT 138.855 0.18 139.115 12.9 ;
      RECT 139.365 0.18 139.625 12.9 ;
      RECT 138.155 136.21 138.355 136.94 ;
      RECT 138.565 136.21 138.925 136.94 ;
      RECT 139.135 136.21 139.335 136.94 ;
      RECT 139.79 136.21 139.99 136.94 ;
      RECT 140.075 0.52 140.335 2.82 ;
      RECT 140.2 136.21 140.56 136.94 ;
      RECT 140.855 136.21 141.055 136.94 ;
      RECT 141.35 136.21 141.71 136.94 ;
      RECT 141.605 0.52 141.865 2.82 ;
      RECT 141.92 136.21 142.12 136.94 ;
      RECT 142.575 136.21 142.775 136.94 ;
      RECT 142.78 0.52 143.04 4.315 ;
      RECT 142.985 136.21 143.345 136.94 ;
      RECT 143.555 136.21 143.755 136.94 ;
      RECT 143.63 0.52 143.89 7.78 ;
      RECT 144.14 0.3 144.4 5.235 ;
      RECT 144.21 136.21 144.41 136.94 ;
      RECT 144.65 0.52 144.91 5.57 ;
      RECT 144.62 136.21 144.98 136.94 ;
      RECT 145.275 136.21 145.475 136.94 ;
      RECT 145.77 136.21 146.13 136.94 ;
      RECT 146.025 0.52 146.285 6.28 ;
      RECT 146.34 136.21 146.54 136.94 ;
      RECT 146.995 136.21 147.195 136.94 ;
      RECT 147.405 136.21 147.765 136.94 ;
      RECT 147.975 136.21 148.175 136.94 ;
      RECT 147.71 0.18 148.48 0.88 ;
      RECT 148.63 136.21 148.83 136.94 ;
      RECT 148.73 0.3 148.99 8.7 ;
      RECT 149.04 136.21 149.4 136.94 ;
      RECT 149.695 136.21 149.895 136.94 ;
      RECT 150.19 136.21 150.55 136.94 ;
      RECT 151.28 0.155 152.05 0.445 ;
      RECT 151.28 0.155 151.54 8.665 ;
      RECT 151.79 0.155 152.05 8.665 ;
      RECT 150.76 136.21 150.96 136.94 ;
      RECT 150.77 0.52 151.03 9.955 ;
      RECT 151.415 136.21 151.615 136.94 ;
      RECT 151.825 136.21 152.185 136.94 ;
      RECT 152.3 0.52 152.56 11.315 ;
      RECT 152.395 136.21 152.595 136.94 ;
      RECT 152.81 0.52 153.07 13.45 ;
      RECT 153.05 136.21 153.25 136.94 ;
      RECT 153.32 0.52 153.58 14.115 ;
      RECT 153.46 136.21 153.82 136.94 ;
      RECT 154.115 136.21 154.315 136.94 ;
      RECT 155.515 0.155 156.285 0.445 ;
      RECT 155.515 0.155 155.775 13.21 ;
      RECT 156.025 0.155 156.285 13.21 ;
      RECT 154.61 136.21 154.97 136.94 ;
      RECT 155.18 136.21 155.38 136.94 ;
      RECT 156.535 0.18 157.305 0.88 ;
      RECT 156.535 0.18 156.795 12.9 ;
      RECT 157.045 0.18 157.305 12.9 ;
      RECT 155.835 136.21 156.035 136.94 ;
      RECT 156.245 136.21 156.605 136.94 ;
      RECT 156.815 136.21 157.015 136.94 ;
      RECT 157.47 136.21 157.67 136.94 ;
      RECT 157.755 0.52 158.015 2.82 ;
      RECT 157.88 136.21 158.24 136.94 ;
      RECT 158.535 136.21 158.735 136.94 ;
      RECT 159.03 136.21 159.39 136.94 ;
      RECT 159.285 0.52 159.545 2.82 ;
      RECT 159.6 136.21 159.8 136.94 ;
      RECT 160.255 136.21 160.455 136.94 ;
      RECT 160.46 0.52 160.72 4.315 ;
      RECT 160.665 136.21 161.025 136.94 ;
      RECT 161.235 136.21 161.435 136.94 ;
      RECT 161.31 0.52 161.57 7.78 ;
      RECT 161.82 0.3 162.08 5.235 ;
      RECT 161.89 136.21 162.09 136.94 ;
      RECT 162.33 0.52 162.59 5.57 ;
      RECT 162.3 136.21 162.66 136.94 ;
      RECT 162.955 136.21 163.155 136.94 ;
      RECT 163.45 136.21 163.81 136.94 ;
      RECT 163.705 0.52 163.965 6.28 ;
      RECT 164.02 136.21 164.22 136.94 ;
      RECT 164.675 136.21 164.875 136.94 ;
      RECT 165.085 136.21 165.445 136.94 ;
      RECT 165.655 136.21 165.855 136.94 ;
      RECT 165.39 0.18 166.16 0.88 ;
      RECT 166.31 136.21 166.51 136.94 ;
      RECT 166.41 0.3 166.67 8.7 ;
      RECT 166.72 136.21 167.08 136.94 ;
      RECT 167.375 136.21 167.575 136.94 ;
      RECT 167.87 136.21 168.23 136.94 ;
      RECT 168.96 0.155 169.73 0.445 ;
      RECT 168.96 0.155 169.22 8.665 ;
      RECT 169.47 0.155 169.73 8.665 ;
      RECT 168.44 136.21 168.64 136.94 ;
      RECT 168.45 0.52 168.71 9.955 ;
      RECT 169.095 136.21 169.295 136.94 ;
      RECT 169.505 136.21 169.865 136.94 ;
      RECT 169.98 0.52 170.24 11.315 ;
      RECT 170.075 136.21 170.275 136.94 ;
      RECT 170.49 0.52 170.75 13.45 ;
      RECT 170.73 136.21 170.93 136.94 ;
      RECT 171 0.52 171.26 14.115 ;
      RECT 171.14 136.21 171.5 136.94 ;
      RECT 171.795 136.21 171.995 136.94 ;
      RECT 173.195 0.155 173.965 0.445 ;
      RECT 173.195 0.155 173.455 13.21 ;
      RECT 173.705 0.155 173.965 13.21 ;
      RECT 172.29 136.21 172.65 136.94 ;
      RECT 172.86 136.21 173.06 136.94 ;
      RECT 174.215 0.18 174.985 0.88 ;
      RECT 174.215 0.18 174.475 12.9 ;
      RECT 174.725 0.18 174.985 12.9 ;
      RECT 173.515 136.21 173.715 136.94 ;
      RECT 173.925 136.21 174.285 136.94 ;
      RECT 174.495 136.21 174.695 136.94 ;
      RECT 175.15 136.21 175.35 136.94 ;
      RECT 175.435 0.52 175.695 2.82 ;
      RECT 175.56 136.21 175.92 136.94 ;
      RECT 176.215 136.21 176.415 136.94 ;
      RECT 176.71 136.21 177.07 136.94 ;
      RECT 176.965 0.52 177.225 2.82 ;
      RECT 177.28 136.21 177.48 136.94 ;
      RECT 177.935 136.21 178.135 136.94 ;
      RECT 178.14 0.52 178.4 4.315 ;
      RECT 178.345 136.21 178.705 136.94 ;
      RECT 178.915 136.21 179.115 136.94 ;
      RECT 178.99 0.52 179.25 7.78 ;
      RECT 179.5 0.3 179.76 5.235 ;
      RECT 179.57 136.21 179.77 136.94 ;
      RECT 180.01 0.52 180.27 5.57 ;
      RECT 179.98 136.21 180.34 136.94 ;
      RECT 180.635 136.21 180.835 136.94 ;
      RECT 181.13 136.21 181.49 136.94 ;
      RECT 181.385 0.52 181.645 6.28 ;
      RECT 181.7 136.21 181.9 136.94 ;
      RECT 182.355 136.21 182.555 136.94 ;
      RECT 182.765 136.21 183.125 136.94 ;
      RECT 183.335 136.21 183.535 136.94 ;
      RECT 183.07 0.18 183.84 0.88 ;
      RECT 183.99 136.21 184.19 136.94 ;
      RECT 184.09 0.3 184.35 8.7 ;
      RECT 184.4 136.21 184.76 136.94 ;
      RECT 185.055 136.21 185.255 136.94 ;
      RECT 185.55 136.21 185.91 136.94 ;
      RECT 186.64 0.155 187.41 0.445 ;
      RECT 186.64 0.155 186.9 8.665 ;
      RECT 187.15 0.155 187.41 8.665 ;
      RECT 186.12 136.21 186.32 136.94 ;
      RECT 186.13 0.52 186.39 9.955 ;
      RECT 186.775 136.21 186.975 136.94 ;
      RECT 187.185 136.21 187.545 136.94 ;
      RECT 187.66 0.52 187.92 11.315 ;
      RECT 187.755 136.21 187.955 136.94 ;
      RECT 188.17 0.52 188.43 13.45 ;
      RECT 188.41 136.21 188.61 136.94 ;
      RECT 188.68 0.52 188.94 14.115 ;
      RECT 188.82 136.21 189.18 136.94 ;
      RECT 189.475 136.21 189.675 136.94 ;
      RECT 190.875 0.155 191.645 0.445 ;
      RECT 190.875 0.155 191.135 13.21 ;
      RECT 191.385 0.155 191.645 13.21 ;
      RECT 189.97 136.21 190.33 136.94 ;
      RECT 190.54 136.21 190.74 136.94 ;
      RECT 191.895 0.18 192.665 0.88 ;
      RECT 191.895 0.18 192.155 12.9 ;
      RECT 192.405 0.18 192.665 12.9 ;
      RECT 191.195 136.21 191.395 136.94 ;
      RECT 191.605 136.21 191.965 136.94 ;
      RECT 192.175 136.21 192.375 136.94 ;
      RECT 192.83 136.21 193.03 136.94 ;
      RECT 193.115 0.52 193.375 2.82 ;
      RECT 193.24 136.21 193.6 136.94 ;
      RECT 193.895 136.21 194.095 136.94 ;
      RECT 194.39 136.21 194.75 136.94 ;
      RECT 194.645 0.52 194.905 2.82 ;
      RECT 194.96 136.21 195.16 136.94 ;
      RECT 195.615 136.21 195.815 136.94 ;
      RECT 195.82 0.52 196.08 4.315 ;
      RECT 196.025 136.21 196.385 136.94 ;
      RECT 196.595 136.21 196.795 136.94 ;
      RECT 196.67 0.52 196.93 7.78 ;
      RECT 197.18 0.3 197.44 5.235 ;
      RECT 197.25 136.21 197.45 136.94 ;
      RECT 197.69 0.52 197.95 5.57 ;
      RECT 197.66 136.21 198.02 136.94 ;
      RECT 198.315 136.21 198.515 136.94 ;
      RECT 198.81 136.21 199.17 136.94 ;
      RECT 199.065 0.52 199.325 6.28 ;
      RECT 199.38 136.21 199.58 136.94 ;
      RECT 200.035 136.21 200.235 136.94 ;
      RECT 200.445 136.21 200.805 136.94 ;
      RECT 201.015 136.21 201.215 136.94 ;
      RECT 200.75 0.18 201.52 0.88 ;
      RECT 201.67 136.21 201.87 136.94 ;
      RECT 201.77 0.3 202.03 8.7 ;
      RECT 202.08 136.21 202.44 136.94 ;
      RECT 202.735 136.21 202.935 136.94 ;
      RECT 203.23 136.21 203.59 136.94 ;
      RECT 204.32 0.155 205.09 0.445 ;
      RECT 204.32 0.155 204.58 8.665 ;
      RECT 204.83 0.155 205.09 8.665 ;
      RECT 203.8 136.21 204 136.94 ;
      RECT 203.81 0.52 204.07 9.955 ;
      RECT 204.455 136.21 204.655 136.94 ;
      RECT 204.865 136.21 205.225 136.94 ;
      RECT 205.34 0.52 205.6 11.315 ;
      RECT 205.435 136.21 205.635 136.94 ;
      RECT 205.85 0.52 206.11 13.45 ;
      RECT 206.09 136.21 206.29 136.94 ;
      RECT 206.36 0.52 206.62 14.115 ;
      RECT 206.5 136.21 206.86 136.94 ;
      RECT 207.155 136.21 207.355 136.94 ;
      RECT 208.555 0.155 209.325 0.445 ;
      RECT 208.555 0.155 208.815 13.21 ;
      RECT 209.065 0.155 209.325 13.21 ;
      RECT 207.65 136.21 208.01 136.94 ;
      RECT 208.22 136.21 208.42 136.94 ;
      RECT 209.575 0.18 210.345 0.88 ;
      RECT 209.575 0.18 209.835 12.9 ;
      RECT 210.085 0.18 210.345 12.9 ;
      RECT 208.875 136.21 209.075 136.94 ;
      RECT 209.285 136.21 209.645 136.94 ;
      RECT 209.855 136.21 210.055 136.94 ;
      RECT 210.51 136.21 210.71 136.94 ;
      RECT 210.795 0.52 211.055 2.82 ;
      RECT 210.92 136.21 211.28 136.94 ;
      RECT 211.575 136.21 211.775 136.94 ;
      RECT 212.07 136.21 212.43 136.94 ;
      RECT 212.325 0.52 212.585 2.82 ;
      RECT 212.64 136.21 212.84 136.94 ;
      RECT 213.295 136.21 213.495 136.94 ;
      RECT 213.5 0.52 213.76 4.315 ;
      RECT 213.705 136.21 214.065 136.94 ;
      RECT 214.275 136.21 214.475 136.94 ;
      RECT 214.35 0.52 214.61 7.78 ;
      RECT 214.86 0.3 215.12 5.235 ;
      RECT 214.93 136.21 215.13 136.94 ;
      RECT 215.37 0.52 215.63 5.57 ;
      RECT 215.34 136.21 215.7 136.94 ;
      RECT 215.995 136.21 216.195 136.94 ;
      RECT 216.49 136.21 216.85 136.94 ;
      RECT 216.745 0.52 217.005 6.28 ;
      RECT 217.06 136.21 217.26 136.94 ;
      RECT 217.715 136.21 217.915 136.94 ;
      RECT 218.125 136.21 218.485 136.94 ;
      RECT 218.695 136.21 218.895 136.94 ;
      RECT 218.43 0.18 219.2 0.88 ;
      RECT 219.35 136.21 219.55 136.94 ;
      RECT 219.45 0.3 219.71 8.7 ;
      RECT 219.76 136.21 220.12 136.94 ;
      RECT 220.415 136.21 220.615 136.94 ;
      RECT 220.91 136.21 221.27 136.94 ;
      RECT 222 0.155 222.77 0.445 ;
      RECT 222 0.155 222.26 8.665 ;
      RECT 222.51 0.155 222.77 8.665 ;
      RECT 221.48 136.21 221.68 136.94 ;
      RECT 221.49 0.52 221.75 9.955 ;
      RECT 222.135 136.21 222.335 136.94 ;
      RECT 222.545 136.21 222.905 136.94 ;
      RECT 223.02 0.52 223.28 11.315 ;
      RECT 223.115 136.21 223.315 136.94 ;
      RECT 223.53 0.52 223.79 13.45 ;
      RECT 223.77 136.21 223.97 136.94 ;
      RECT 224.04 0.52 224.3 14.115 ;
      RECT 224.18 136.21 224.54 136.94 ;
      RECT 224.835 136.21 225.035 136.94 ;
      RECT 226.235 0.155 227.005 0.445 ;
      RECT 226.235 0.155 226.495 13.21 ;
      RECT 226.745 0.155 227.005 13.21 ;
      RECT 225.33 136.21 225.69 136.94 ;
      RECT 225.9 136.21 226.1 136.94 ;
      RECT 227.255 0.18 228.025 0.88 ;
      RECT 227.255 0.18 227.515 12.9 ;
      RECT 227.765 0.18 228.025 12.9 ;
      RECT 226.555 136.21 226.755 136.94 ;
      RECT 226.965 136.21 227.325 136.94 ;
      RECT 227.535 136.21 227.735 136.94 ;
      RECT 228.19 136.21 228.39 136.94 ;
      RECT 228.475 0.52 228.735 2.82 ;
      RECT 228.6 136.21 228.96 136.94 ;
      RECT 229.255 136.21 229.455 136.94 ;
      RECT 229.75 136.21 230.11 136.94 ;
      RECT 230.005 0.52 230.265 2.82 ;
      RECT 230.32 136.21 230.52 136.94 ;
      RECT 230.975 136.21 231.175 136.94 ;
      RECT 231.18 0.52 231.44 4.315 ;
      RECT 231.385 136.21 231.745 136.94 ;
      RECT 231.955 136.21 232.155 136.94 ;
      RECT 232.03 0.52 232.29 7.78 ;
      RECT 232.54 0.3 232.8 5.235 ;
      RECT 232.61 136.21 232.81 136.94 ;
      RECT 233.05 0.52 233.31 5.57 ;
      RECT 233.02 136.21 233.38 136.94 ;
      RECT 233.675 136.21 233.875 136.94 ;
      RECT 234.17 136.21 234.53 136.94 ;
      RECT 234.425 0.52 234.685 6.28 ;
      RECT 234.74 136.21 234.94 136.94 ;
      RECT 235.395 136.21 235.595 136.94 ;
      RECT 235.805 136.21 236.165 136.94 ;
      RECT 236.375 136.21 236.575 136.94 ;
      RECT 236.11 0.18 236.88 0.88 ;
      RECT 237.03 136.21 237.23 136.94 ;
      RECT 237.13 0.3 237.39 8.7 ;
      RECT 237.44 136.21 237.8 136.94 ;
      RECT 238.095 136.21 238.295 136.94 ;
      RECT 238.59 136.21 238.95 136.94 ;
      RECT 239.68 0.155 240.45 0.445 ;
      RECT 239.68 0.155 239.94 8.665 ;
      RECT 240.19 0.155 240.45 8.665 ;
      RECT 239.16 136.21 239.36 136.94 ;
      RECT 239.17 0.52 239.43 9.955 ;
      RECT 239.815 136.21 240.015 136.94 ;
      RECT 240.225 136.21 240.585 136.94 ;
      RECT 240.7 0.52 240.96 11.315 ;
      RECT 240.795 136.21 240.995 136.94 ;
      RECT 241.21 0.52 241.47 13.45 ;
      RECT 241.45 136.21 241.65 136.94 ;
      RECT 241.72 0.52 241.98 14.115 ;
      RECT 241.86 136.21 242.22 136.94 ;
      RECT 242.515 136.21 242.715 136.94 ;
      RECT 243.915 0.155 244.685 0.445 ;
      RECT 243.915 0.155 244.175 13.21 ;
      RECT 244.425 0.155 244.685 13.21 ;
      RECT 243.01 136.21 243.37 136.94 ;
      RECT 243.58 136.21 243.78 136.94 ;
      RECT 244.935 0.18 245.705 0.88 ;
      RECT 244.935 0.18 245.195 12.9 ;
      RECT 245.445 0.18 245.705 12.9 ;
      RECT 244.235 136.21 244.435 136.94 ;
      RECT 244.645 136.21 245.005 136.94 ;
      RECT 245.215 136.21 245.415 136.94 ;
      RECT 245.87 136.21 246.07 136.94 ;
      RECT 246.155 0.52 246.415 2.82 ;
      RECT 246.28 136.21 246.64 136.94 ;
      RECT 246.935 136.21 247.135 136.94 ;
      RECT 247.43 136.21 247.79 136.94 ;
      RECT 247.685 0.52 247.945 2.82 ;
      RECT 248 136.21 248.2 136.94 ;
      RECT 248.655 136.21 248.855 136.94 ;
      RECT 248.86 0.52 249.12 4.315 ;
      RECT 249.065 136.21 249.425 136.94 ;
      RECT 249.635 136.21 249.835 136.94 ;
      RECT 249.71 0.52 249.97 7.78 ;
      RECT 250.22 0.3 250.48 5.235 ;
      RECT 250.29 136.21 250.49 136.94 ;
      RECT 250.73 0.52 250.99 5.57 ;
      RECT 250.7 136.21 251.06 136.94 ;
      RECT 251.355 136.21 251.555 136.94 ;
      RECT 251.85 136.21 252.21 136.94 ;
      RECT 252.105 0.52 252.365 6.28 ;
      RECT 252.42 136.21 252.62 136.94 ;
      RECT 253.075 136.21 253.275 136.94 ;
      RECT 253.485 136.21 253.845 136.94 ;
      RECT 254.055 136.21 254.255 136.94 ;
      RECT 253.79 0.18 254.56 0.88 ;
      RECT 254.71 136.21 254.91 136.94 ;
      RECT 254.81 0.3 255.07 8.7 ;
      RECT 255.12 136.21 255.48 136.94 ;
      RECT 255.775 136.21 255.975 136.94 ;
      RECT 256.27 136.21 256.63 136.94 ;
      RECT 257.36 0.155 258.13 0.445 ;
      RECT 257.36 0.155 257.62 8.665 ;
      RECT 257.87 0.155 258.13 8.665 ;
      RECT 256.84 136.21 257.04 136.94 ;
      RECT 256.85 0.52 257.11 9.955 ;
      RECT 257.495 136.21 257.695 136.94 ;
      RECT 257.905 136.21 258.265 136.94 ;
      RECT 258.38 0.52 258.64 11.315 ;
      RECT 258.475 136.21 258.675 136.94 ;
      RECT 258.89 0.52 259.15 13.45 ;
      RECT 259.13 136.21 259.33 136.94 ;
      RECT 259.4 0.52 259.66 14.115 ;
      RECT 259.54 136.21 259.9 136.94 ;
      RECT 260.195 136.21 260.395 136.94 ;
      RECT 261.595 0.155 262.365 0.445 ;
      RECT 261.595 0.155 261.855 13.21 ;
      RECT 262.105 0.155 262.365 13.21 ;
      RECT 260.69 136.21 261.05 136.94 ;
      RECT 261.26 136.21 261.46 136.94 ;
      RECT 262.615 0.18 263.385 0.88 ;
      RECT 262.615 0.18 262.875 12.9 ;
      RECT 263.125 0.18 263.385 12.9 ;
      RECT 261.915 136.21 262.115 136.94 ;
      RECT 262.325 136.21 262.685 136.94 ;
      RECT 262.895 136.21 263.095 136.94 ;
      RECT 263.55 136.21 263.75 136.94 ;
      RECT 263.835 0.52 264.095 2.82 ;
      RECT 263.96 136.21 264.32 136.94 ;
      RECT 264.615 136.21 264.815 136.94 ;
      RECT 265.11 136.21 265.47 136.94 ;
      RECT 265.365 0.52 265.625 2.82 ;
      RECT 265.68 136.21 265.88 136.94 ;
      RECT 266.335 136.21 266.535 136.94 ;
      RECT 266.54 0.52 266.8 4.315 ;
      RECT 266.745 136.21 267.105 136.94 ;
      RECT 267.315 136.21 267.515 136.94 ;
      RECT 267.39 0.52 267.65 7.78 ;
      RECT 267.9 0.3 268.16 5.235 ;
      RECT 267.97 136.21 268.17 136.94 ;
      RECT 268.41 0.52 268.67 5.57 ;
      RECT 268.38 136.21 268.74 136.94 ;
      RECT 269.035 136.21 269.235 136.94 ;
      RECT 269.53 136.21 269.89 136.94 ;
      RECT 269.785 0.52 270.045 6.28 ;
      RECT 270.1 136.21 270.3 136.94 ;
      RECT 270.755 136.21 270.955 136.94 ;
      RECT 271.165 136.21 271.525 136.94 ;
      RECT 271.735 136.21 271.935 136.94 ;
      RECT 271.47 0.18 272.24 0.88 ;
      RECT 272.39 136.21 272.59 136.94 ;
      RECT 272.49 0.3 272.75 8.7 ;
      RECT 272.8 136.21 273.16 136.94 ;
      RECT 273.455 136.21 273.655 136.94 ;
      RECT 273.95 136.21 274.31 136.94 ;
      RECT 275.04 0.155 275.81 0.445 ;
      RECT 275.04 0.155 275.3 8.665 ;
      RECT 275.55 0.155 275.81 8.665 ;
      RECT 274.52 136.21 274.72 136.94 ;
      RECT 274.53 0.52 274.79 9.955 ;
      RECT 275.175 136.21 275.375 136.94 ;
      RECT 275.585 136.21 275.945 136.94 ;
      RECT 276.06 0.52 276.32 11.315 ;
      RECT 276.155 136.21 276.355 136.94 ;
      RECT 276.57 0.52 276.83 13.45 ;
      RECT 276.81 136.21 277.01 136.94 ;
      RECT 277.08 0.52 277.34 14.115 ;
      RECT 277.22 136.21 277.58 136.94 ;
      RECT 277.875 136.21 278.075 136.94 ;
      RECT 279.275 0.155 280.045 0.445 ;
      RECT 279.275 0.155 279.535 13.21 ;
      RECT 279.785 0.155 280.045 13.21 ;
      RECT 278.37 136.21 278.73 136.94 ;
      RECT 278.94 136.21 279.14 136.94 ;
      RECT 280.295 0.18 281.065 0.88 ;
      RECT 280.295 0.18 280.555 12.9 ;
      RECT 280.805 0.18 281.065 12.9 ;
      RECT 279.595 136.21 279.795 136.94 ;
      RECT 280.005 136.21 280.365 136.94 ;
      RECT 280.575 136.21 280.775 136.94 ;
      RECT 281.23 136.21 281.43 136.94 ;
      RECT 281.515 0.52 281.775 2.82 ;
      RECT 281.64 136.21 282 136.94 ;
      RECT 282.295 136.21 282.495 136.94 ;
      RECT 282.79 136.21 283.15 136.94 ;
      RECT 283.045 0.52 283.305 2.82 ;
      RECT 283.36 136.21 283.56 136.94 ;
      RECT 284.015 136.21 284.215 136.94 ;
      RECT 284.22 0.52 284.48 4.315 ;
      RECT 285.75 0.17 286.52 0.43 ;
      RECT 285.75 0.17 286.01 8.7 ;
      RECT 286.26 0.17 286.52 8.7 ;
      RECT 286.77 0.18 287.54 0.88 ;
      RECT 286.77 0.18 287.03 8.7 ;
      RECT 287.28 0.18 287.54 8.7 ;
      RECT 287.79 0.17 288.56 0.43 ;
      RECT 287.79 0.17 288.05 8.7 ;
      RECT 288.3 0.17 288.56 8.7 ;
      RECT 288.81 0.18 289.58 0.88 ;
      RECT 288.81 0.18 289.07 8.7 ;
      RECT 289.32 0.18 289.58 8.7 ;
      RECT 289.83 0.17 290.6 0.43 ;
      RECT 289.83 0.17 290.09 8.7 ;
      RECT 290.34 0.17 290.6 8.7 ;
      RECT 290.85 0.18 291.62 0.88 ;
      RECT 290.85 0.18 291.11 8.7 ;
      RECT 291.36 0.18 291.62 8.7 ;
      RECT 291.87 0.17 292.64 0.43 ;
      RECT 291.87 0.17 292.13 8.7 ;
      RECT 292.38 0.17 292.64 8.7 ;
      RECT 292.89 0.18 293.66 0.88 ;
      RECT 292.89 0.18 293.15 8.7 ;
      RECT 293.4 0.18 293.66 8.7 ;
      RECT 293.91 0.17 294.68 0.43 ;
      RECT 293.91 0.17 294.17 8.7 ;
      RECT 294.42 0.17 294.68 8.7 ;
      RECT 294.93 0.18 295.7 0.88 ;
      RECT 294.93 0.18 295.19 8.7 ;
      RECT 295.44 0.18 295.7 8.7 ;
      RECT 295.95 0.17 296.72 0.43 ;
      RECT 295.95 0.17 296.21 8.7 ;
      RECT 296.46 0.17 296.72 8.7 ;
      RECT 296.97 0.18 297.74 0.88 ;
      RECT 296.97 0.18 297.23 8.7 ;
      RECT 297.48 0.18 297.74 8.7 ;
      RECT 297.99 0.17 298.76 0.43 ;
      RECT 297.99 0.17 298.25 8.7 ;
      RECT 298.5 0.17 298.76 8.7 ;
      RECT 299.01 0.18 299.78 0.88 ;
      RECT 299.01 0.18 299.27 8.7 ;
      RECT 299.52 0.18 299.78 8.7 ;
      RECT 300.03 0.17 300.8 0.43 ;
      RECT 300.03 0.17 300.29 8.7 ;
      RECT 300.54 0.17 300.8 8.7 ;
      RECT 301.05 0.18 301.82 0.88 ;
      RECT 301.05 0.18 301.31 8.7 ;
      RECT 301.56 0.18 301.82 8.7 ;
      RECT 302.07 0.17 302.84 0.43 ;
      RECT 302.07 0.17 302.33 8.7 ;
      RECT 302.58 0.17 302.84 8.7 ;
      RECT 303.09 0.18 303.86 0.88 ;
      RECT 303.09 0.18 303.35 8.7 ;
      RECT 303.6 0.18 303.86 8.7 ;
      RECT 304.11 0.17 304.88 0.43 ;
      RECT 304.11 0.17 304.37 8.7 ;
      RECT 304.62 0.17 304.88 8.7 ;
      RECT 305.13 0.18 305.9 0.88 ;
      RECT 305.13 0.18 305.39 8.7 ;
      RECT 305.64 0.18 305.9 8.7 ;
      RECT 306.15 0.17 306.92 0.43 ;
      RECT 306.15 0.17 306.41 8.7 ;
      RECT 306.66 0.17 306.92 8.7 ;
      RECT 307.17 0.18 307.94 0.88 ;
      RECT 307.17 0.18 307.43 8.7 ;
      RECT 307.68 0.18 307.94 8.7 ;
      RECT 308.19 0.17 308.96 0.43 ;
      RECT 308.19 0.17 308.45 8.7 ;
      RECT 308.7 0.17 308.96 8.7 ;
      RECT 309.21 0.18 309.98 0.88 ;
      RECT 309.21 0.18 309.47 8.7 ;
      RECT 309.72 0.18 309.98 8.7 ;
      RECT 284.425 136.21 284.785 136.94 ;
      RECT 284.995 136.21 285.195 136.94 ;
      RECT 311.605 0.18 312.375 0.88 ;
      RECT 311.605 0.18 311.865 8.7 ;
      RECT 312.115 0.18 312.375 8.7 ;
      RECT 312.625 0.17 313.395 0.43 ;
      RECT 312.625 0.17 312.885 8.7 ;
      RECT 313.135 0.17 313.395 8.7 ;
      RECT 285.82 136.13 286.02 136.94 ;
      RECT 310.585 0.3 310.845 8.7 ;
      RECT 314.665 0.18 315.435 0.88 ;
      RECT 314.665 0.18 314.925 8.7 ;
      RECT 315.175 0.18 315.435 8.7 ;
      RECT 311.095 0.3 311.355 8.7 ;
      RECT 313.645 0 313.905 8.7 ;
      RECT 314.155 0 314.415 8.7 ;
      RECT 315.685 0.52 315.945 8.7 ;
      RECT 316.195 0.3 316.455 8.7 ;
      RECT 316.705 0.3 316.965 8.7 ;
      RECT 317.215 0.3 317.475 8.7 ;
      RECT 317.725 0.3 317.985 8.7 ;
      RECT 318.235 0.3 318.495 8.7 ;
      RECT 318.745 0.3 319.005 8.7 ;
      RECT 319.255 0.3 319.515 8.7 ;
      RECT 321.295 0.18 322.065 0.88 ;
      RECT 321.295 0.18 321.555 8.7 ;
      RECT 321.805 0.18 322.065 8.7 ;
      RECT 319.765 0.3 320.025 8.7 ;
      RECT 320.275 0 320.535 8.7 ;
      RECT 320.785 0 321.045 8.7 ;
      RECT 322.315 0 322.575 8.7 ;
      RECT 322.825 0 323.085 8.7 ;
      RECT 323.335 0.52 323.595 8.7 ;
      RECT 323.845 0.52 324.105 8.7 ;
      RECT 324.355 0.52 324.615 8.7 ;
      RECT 324.865 0.52 325.125 8.7 ;
      RECT 325.375 0.52 325.635 8.7 ;
      RECT 325.885 0.52 326.145 8.7 ;
      RECT 326.395 0.52 326.655 8.7 ;
      RECT 326.905 0.52 327.165 8.7 ;
      RECT 327.415 0.3 327.675 8.7 ;
      RECT 327.925 0.3 328.185 8.7 ;
      RECT 328.435 0.3 328.695 8.7 ;
      RECT 328.945 0.52 329.205 8.7 ;
      RECT 329.455 0.52 329.715 8.7 ;
      RECT 329.965 0.3 330.225 8.7 ;
      RECT 330.475 0.3 330.735 8.7 ;
      RECT 330.985 0.3 331.245 8.7 ;
      RECT 331.495 0.52 331.755 8.7 ;
      RECT 332.005 0.52 332.265 8.7 ;
      RECT 332.515 0.3 332.775 8.7 ;
      RECT 333.025 0.52 333.285 8.7 ;
      RECT 333.535 0.52 333.795 8.7 ;
      RECT 334.045 0.52 334.305 8.7 ;
      RECT 334.555 0.52 334.815 8.7 ;
      RECT 335.065 0.52 335.325 8.7 ;
      RECT 335.575 0.3 335.835 8.7 ;
      RECT 336.085 0.52 336.345 8.7 ;
      RECT 336.595 0.52 336.855 8.7 ;
      RECT 337.105 0.3 337.365 8.7 ;
      RECT 337.615 0.52 337.875 8.7 ;
      RECT 339.655 0.17 340.425 0.43 ;
      RECT 339.655 0.17 339.915 8.7 ;
      RECT 340.165 0.17 340.425 8.7 ;
      RECT 338.125 0.52 338.385 8.7 ;
      RECT 338.635 0.3 338.895 8.7 ;
      RECT 339.145 0.3 339.405 8.7 ;
      RECT 342.205 0.17 342.975 0.43 ;
      RECT 342.205 0.17 342.465 8.7 ;
      RECT 342.715 0.17 342.975 8.7 ;
      RECT 340.675 0.3 340.935 8.7 ;
      RECT 343.735 0.18 344.505 0.88 ;
      RECT 343.735 0.18 343.995 8.7 ;
      RECT 344.245 0.18 344.505 8.7 ;
      RECT 341.185 0.3 341.445 8.7 ;
      RECT 341.695 0.3 341.955 8.7 ;
      RECT 343.225 0.3 343.485 8.7 ;
      RECT 344.755 0 345.015 8.7 ;
      RECT 345.265 0 345.525 8.7 ;
      RECT 345.775 0.52 346.035 8.7 ;
      RECT 346.285 0.52 346.545 8.7 ;
      RECT 346.795 0.52 347.055 8.7 ;
      RECT 347.305 0.52 347.565 8.7 ;
      RECT 347.815 0 348.075 8.7 ;
      RECT 348.325 0 348.585 8.7 ;
      RECT 348.835 0.3 349.095 8.7 ;
      RECT 349.345 0.3 349.605 8.7 ;
      RECT 349.855 0 350.115 8.7 ;
      RECT 350.365 0 350.625 8.7 ;
      RECT 350.875 0.3 351.135 8.7 ;
      RECT 351.695 0.3 351.955 8.7 ;
      RECT 352.205 0 352.465 8.7 ;
      RECT 352.715 0 352.975 8.7 ;
      RECT 353.225 0.3 353.485 8.7 ;
      RECT 353.735 0.3 353.995 8.7 ;
      RECT 354.245 0 354.505 8.7 ;
      RECT 354.755 0 355.015 8.7 ;
      RECT 355.265 0.52 355.525 8.7 ;
      RECT 355.775 0.52 356.035 8.7 ;
      RECT 356.285 0.52 356.545 8.7 ;
      RECT 358.325 0.18 359.095 0.88 ;
      RECT 358.325 0.18 358.585 8.7 ;
      RECT 358.835 0.18 359.095 8.7 ;
      RECT 356.795 0.52 357.055 8.7 ;
      RECT 359.855 0.17 360.625 0.43 ;
      RECT 359.855 0.17 360.115 8.7 ;
      RECT 360.365 0.17 360.625 8.7 ;
      RECT 357.305 0 357.565 8.7 ;
      RECT 357.815 0 358.075 8.7 ;
      RECT 359.345 0.3 359.605 8.7 ;
      RECT 362.405 0.17 363.175 0.43 ;
      RECT 362.405 0.17 362.665 8.7 ;
      RECT 362.915 0.17 363.175 8.7 ;
      RECT 360.875 0.3 361.135 8.7 ;
      RECT 361.385 0.3 361.645 8.7 ;
      RECT 361.895 0.3 362.155 8.7 ;
      RECT 363.425 0.3 363.685 8.7 ;
      RECT 363.935 0.3 364.195 8.7 ;
      RECT 364.445 0.52 364.705 8.7 ;
      RECT 364.955 0.52 365.215 8.7 ;
      RECT 365.465 0.3 365.725 8.7 ;
      RECT 365.975 0.52 366.235 8.7 ;
      RECT 366.485 0.52 366.745 8.7 ;
      RECT 366.995 0.3 367.255 8.7 ;
      RECT 367.505 0.52 367.765 8.7 ;
      RECT 368.015 0.52 368.275 8.7 ;
      RECT 368.525 0.52 368.785 8.7 ;
      RECT 369.035 0.52 369.295 8.7 ;
      RECT 369.545 0.52 369.805 8.7 ;
      RECT 370.055 0.3 370.315 8.7 ;
      RECT 370.565 0.52 370.825 8.7 ;
      RECT 371.075 0.52 371.335 8.7 ;
      RECT 371.585 0.3 371.845 8.7 ;
      RECT 372.095 0.3 372.355 8.7 ;
      RECT 372.605 0.3 372.865 8.7 ;
      RECT 373.115 0.52 373.375 8.7 ;
      RECT 373.625 0.52 373.885 8.7 ;
      RECT 374.135 0.3 374.395 8.7 ;
      RECT 374.645 0.3 374.905 8.7 ;
      RECT 375.155 0.3 375.415 8.7 ;
      RECT 375.665 0.52 375.925 8.7 ;
      RECT 376.175 0.52 376.435 8.7 ;
      RECT 376.685 0.52 376.945 8.7 ;
      RECT 377.195 0.52 377.455 8.7 ;
      RECT 377.705 0.52 377.965 8.7 ;
      RECT 378.215 0.52 378.475 8.7 ;
      RECT 378.725 0.52 378.985 8.7 ;
      RECT 380.765 0.18 381.535 0.88 ;
      RECT 380.765 0.18 381.025 8.7 ;
      RECT 381.275 0.18 381.535 8.7 ;
      RECT 379.235 0.52 379.495 8.7 ;
      RECT 379.745 0 380.005 8.7 ;
      RECT 380.255 0 380.515 8.7 ;
      RECT 381.785 0 382.045 8.7 ;
      RECT 382.295 0 382.555 8.7 ;
      RECT 382.805 0.3 383.065 8.7 ;
      RECT 383.315 0.3 383.575 8.7 ;
      RECT 383.825 0.3 384.085 8.7 ;
      RECT 384.335 0.3 384.595 8.7 ;
      RECT 384.845 0.3 385.105 8.7 ;
      RECT 385.355 0.3 385.615 8.7 ;
      RECT 387.395 0.18 388.165 0.88 ;
      RECT 387.395 0.18 387.655 8.7 ;
      RECT 387.905 0.18 388.165 8.7 ;
      RECT 385.865 0.3 386.125 8.7 ;
      RECT 386.375 0.3 386.635 8.7 ;
      RECT 389.435 0.17 390.205 0.43 ;
      RECT 389.435 0.17 389.695 8.7 ;
      RECT 389.945 0.17 390.205 8.7 ;
      RECT 390.455 0.18 391.225 0.88 ;
      RECT 390.455 0.18 390.715 8.7 ;
      RECT 390.965 0.18 391.225 8.7 ;
      RECT 386.885 0.52 387.145 8.7 ;
      RECT 388.415 0 388.675 8.7 ;
      RECT 392.85 0.18 393.62 0.88 ;
      RECT 392.85 0.18 393.11 8.7 ;
      RECT 393.36 0.18 393.62 8.7 ;
      RECT 393.87 0.17 394.64 0.43 ;
      RECT 393.87 0.17 394.13 8.7 ;
      RECT 394.38 0.17 394.64 8.7 ;
      RECT 394.89 0.18 395.66 0.88 ;
      RECT 394.89 0.18 395.15 8.7 ;
      RECT 395.4 0.18 395.66 8.7 ;
      RECT 395.91 0.17 396.68 0.43 ;
      RECT 395.91 0.17 396.17 8.7 ;
      RECT 396.42 0.17 396.68 8.7 ;
      RECT 396.93 0.18 397.7 0.88 ;
      RECT 396.93 0.18 397.19 8.7 ;
      RECT 397.44 0.18 397.7 8.7 ;
      RECT 397.95 0.17 398.72 0.43 ;
      RECT 397.95 0.17 398.21 8.7 ;
      RECT 398.46 0.17 398.72 8.7 ;
      RECT 398.97 0.18 399.74 0.88 ;
      RECT 398.97 0.18 399.23 8.7 ;
      RECT 399.48 0.18 399.74 8.7 ;
      RECT 399.99 0.17 400.76 0.43 ;
      RECT 399.99 0.17 400.25 8.7 ;
      RECT 400.5 0.17 400.76 8.7 ;
      RECT 401.01 0.18 401.78 0.88 ;
      RECT 401.01 0.18 401.27 8.7 ;
      RECT 401.52 0.18 401.78 8.7 ;
      RECT 402.03 0.17 402.8 0.43 ;
      RECT 402.03 0.17 402.29 8.7 ;
      RECT 402.54 0.17 402.8 8.7 ;
      RECT 403.05 0.18 403.82 0.88 ;
      RECT 403.05 0.18 403.31 8.7 ;
      RECT 403.56 0.18 403.82 8.7 ;
      RECT 404.07 0.17 404.84 0.43 ;
      RECT 404.07 0.17 404.33 8.7 ;
      RECT 404.58 0.17 404.84 8.7 ;
      RECT 405.09 0.18 405.86 0.88 ;
      RECT 405.09 0.18 405.35 8.7 ;
      RECT 405.6 0.18 405.86 8.7 ;
      RECT 406.11 0.17 406.88 0.43 ;
      RECT 406.11 0.17 406.37 8.7 ;
      RECT 406.62 0.17 406.88 8.7 ;
      RECT 407.13 0.18 407.9 0.88 ;
      RECT 407.13 0.18 407.39 8.7 ;
      RECT 407.64 0.18 407.9 8.7 ;
      RECT 408.15 0.17 408.92 0.43 ;
      RECT 408.15 0.17 408.41 8.7 ;
      RECT 408.66 0.17 408.92 8.7 ;
      RECT 409.17 0.18 409.94 0.88 ;
      RECT 409.17 0.18 409.43 8.7 ;
      RECT 409.68 0.18 409.94 8.7 ;
      RECT 410.19 0.17 410.96 0.43 ;
      RECT 410.19 0.17 410.45 8.7 ;
      RECT 410.7 0.17 410.96 8.7 ;
      RECT 411.21 0.18 411.98 0.88 ;
      RECT 411.21 0.18 411.47 8.7 ;
      RECT 411.72 0.18 411.98 8.7 ;
      RECT 412.23 0.17 413 0.43 ;
      RECT 412.23 0.17 412.49 8.7 ;
      RECT 412.74 0.17 413 8.7 ;
      RECT 413.25 0.18 414.02 0.88 ;
      RECT 413.25 0.18 413.51 8.7 ;
      RECT 413.76 0.18 414.02 8.7 ;
      RECT 414.27 0.17 415.04 0.43 ;
      RECT 414.27 0.17 414.53 8.7 ;
      RECT 414.78 0.17 415.04 8.7 ;
      RECT 415.29 0.18 416.06 0.88 ;
      RECT 415.29 0.18 415.55 8.7 ;
      RECT 415.8 0.18 416.06 8.7 ;
      RECT 388.925 0 389.185 8.7 ;
      RECT 416.31 0.17 417.08 0.43 ;
      RECT 416.31 0.17 416.57 8.7 ;
      RECT 416.82 0.17 417.08 8.7 ;
      RECT 391.475 0.3 391.735 8.7 ;
      RECT 391.985 0.3 392.245 8.7 ;
      RECT 416.81 136.13 417.01 136.94 ;
      RECT 417.635 136.21 417.835 136.94 ;
      RECT 418.045 136.21 418.405 136.94 ;
      RECT 418.35 0.52 418.61 4.315 ;
      RECT 418.615 136.21 418.815 136.94 ;
      RECT 419.27 136.21 419.47 136.94 ;
      RECT 419.525 0.52 419.785 2.82 ;
      RECT 419.68 136.21 420.04 136.94 ;
      RECT 420.335 136.21 420.535 136.94 ;
      RECT 420.83 136.21 421.19 136.94 ;
      RECT 421.765 0.18 422.535 0.88 ;
      RECT 421.765 0.18 422.025 12.9 ;
      RECT 422.275 0.18 422.535 12.9 ;
      RECT 421.055 0.52 421.315 2.82 ;
      RECT 421.4 136.21 421.6 136.94 ;
      RECT 422.785 0.155 423.555 0.445 ;
      RECT 422.785 0.155 423.045 13.21 ;
      RECT 423.295 0.155 423.555 13.21 ;
      RECT 422.055 136.21 422.255 136.94 ;
      RECT 422.465 136.21 422.825 136.94 ;
      RECT 423.035 136.21 423.235 136.94 ;
      RECT 423.69 136.21 423.89 136.94 ;
      RECT 424.1 136.21 424.46 136.94 ;
      RECT 424.755 136.21 424.955 136.94 ;
      RECT 425.25 136.21 425.61 136.94 ;
      RECT 425.49 0.52 425.75 14.115 ;
      RECT 425.82 136.21 426.02 136.94 ;
      RECT 426 0.52 426.26 13.45 ;
      RECT 426.475 136.21 426.675 136.94 ;
      RECT 427.02 0.155 427.79 0.445 ;
      RECT 427.02 0.155 427.28 8.665 ;
      RECT 427.53 0.155 427.79 8.665 ;
      RECT 426.51 0.52 426.77 11.315 ;
      RECT 426.885 136.21 427.245 136.94 ;
      RECT 427.455 136.21 427.655 136.94 ;
      RECT 428.04 0.52 428.3 9.955 ;
      RECT 428.11 136.21 428.31 136.94 ;
      RECT 428.52 136.21 428.88 136.94 ;
      RECT 429.175 136.21 429.375 136.94 ;
      RECT 429.67 136.21 430.03 136.94 ;
      RECT 430.08 0.3 430.34 8.7 ;
      RECT 430.24 136.21 430.44 136.94 ;
      RECT 430.895 136.21 431.095 136.94 ;
      RECT 430.59 0.18 431.36 0.88 ;
      RECT 431.305 136.21 431.665 136.94 ;
      RECT 431.875 136.21 432.075 136.94 ;
      RECT 432.53 136.21 432.73 136.94 ;
      RECT 432.785 0.52 433.045 6.28 ;
      RECT 432.94 136.21 433.3 136.94 ;
      RECT 433.595 136.21 433.795 136.94 ;
      RECT 434.16 0.52 434.42 5.57 ;
      RECT 434.09 136.21 434.45 136.94 ;
      RECT 434.66 136.21 434.86 136.94 ;
      RECT 434.67 0.3 434.93 5.235 ;
      RECT 435.18 0.52 435.44 7.78 ;
      RECT 435.315 136.21 435.515 136.94 ;
      RECT 435.725 136.21 436.085 136.94 ;
      RECT 436.03 0.52 436.29 4.315 ;
      RECT 436.295 136.21 436.495 136.94 ;
      RECT 436.95 136.21 437.15 136.94 ;
      RECT 437.205 0.52 437.465 2.82 ;
      RECT 437.36 136.21 437.72 136.94 ;
      RECT 438.015 136.21 438.215 136.94 ;
      RECT 438.51 136.21 438.87 136.94 ;
      RECT 439.445 0.18 440.215 0.88 ;
      RECT 439.445 0.18 439.705 12.9 ;
      RECT 439.955 0.18 440.215 12.9 ;
      RECT 438.735 0.52 438.995 2.82 ;
      RECT 439.08 136.21 439.28 136.94 ;
      RECT 440.465 0.155 441.235 0.445 ;
      RECT 440.465 0.155 440.725 13.21 ;
      RECT 440.975 0.155 441.235 13.21 ;
      RECT 439.735 136.21 439.935 136.94 ;
      RECT 440.145 136.21 440.505 136.94 ;
      RECT 440.715 136.21 440.915 136.94 ;
      RECT 441.37 136.21 441.57 136.94 ;
      RECT 441.78 136.21 442.14 136.94 ;
      RECT 442.435 136.21 442.635 136.94 ;
      RECT 442.93 136.21 443.29 136.94 ;
      RECT 443.17 0.52 443.43 14.115 ;
      RECT 443.5 136.21 443.7 136.94 ;
      RECT 443.68 0.52 443.94 13.45 ;
      RECT 444.155 136.21 444.355 136.94 ;
      RECT 444.7 0.155 445.47 0.445 ;
      RECT 444.7 0.155 444.96 8.665 ;
      RECT 445.21 0.155 445.47 8.665 ;
      RECT 444.19 0.52 444.45 11.315 ;
      RECT 444.565 136.21 444.925 136.94 ;
      RECT 445.135 136.21 445.335 136.94 ;
      RECT 445.72 0.52 445.98 9.955 ;
      RECT 445.79 136.21 445.99 136.94 ;
      RECT 446.2 136.21 446.56 136.94 ;
      RECT 446.855 136.21 447.055 136.94 ;
      RECT 447.35 136.21 447.71 136.94 ;
      RECT 447.76 0.3 448.02 8.7 ;
      RECT 447.92 136.21 448.12 136.94 ;
      RECT 448.575 136.21 448.775 136.94 ;
      RECT 448.27 0.18 449.04 0.88 ;
      RECT 448.985 136.21 449.345 136.94 ;
      RECT 449.555 136.21 449.755 136.94 ;
      RECT 450.21 136.21 450.41 136.94 ;
      RECT 450.465 0.52 450.725 6.28 ;
      RECT 450.62 136.21 450.98 136.94 ;
      RECT 451.275 136.21 451.475 136.94 ;
      RECT 451.84 0.52 452.1 5.57 ;
      RECT 451.77 136.21 452.13 136.94 ;
      RECT 452.34 136.21 452.54 136.94 ;
      RECT 452.35 0.3 452.61 5.235 ;
      RECT 452.86 0.52 453.12 7.78 ;
      RECT 452.995 136.21 453.195 136.94 ;
      RECT 453.405 136.21 453.765 136.94 ;
      RECT 453.71 0.52 453.97 4.315 ;
      RECT 453.975 136.21 454.175 136.94 ;
      RECT 454.63 136.21 454.83 136.94 ;
      RECT 454.885 0.52 455.145 2.82 ;
      RECT 455.04 136.21 455.4 136.94 ;
      RECT 455.695 136.21 455.895 136.94 ;
      RECT 456.19 136.21 456.55 136.94 ;
      RECT 457.125 0.18 457.895 0.88 ;
      RECT 457.125 0.18 457.385 12.9 ;
      RECT 457.635 0.18 457.895 12.9 ;
      RECT 456.415 0.52 456.675 2.82 ;
      RECT 456.76 136.21 456.96 136.94 ;
      RECT 458.145 0.155 458.915 0.445 ;
      RECT 458.145 0.155 458.405 13.21 ;
      RECT 458.655 0.155 458.915 13.21 ;
      RECT 457.415 136.21 457.615 136.94 ;
      RECT 457.825 136.21 458.185 136.94 ;
      RECT 458.395 136.21 458.595 136.94 ;
      RECT 459.05 136.21 459.25 136.94 ;
      RECT 459.46 136.21 459.82 136.94 ;
      RECT 460.115 136.21 460.315 136.94 ;
      RECT 460.61 136.21 460.97 136.94 ;
      RECT 460.85 0.52 461.11 14.115 ;
      RECT 461.18 136.21 461.38 136.94 ;
      RECT 461.36 0.52 461.62 13.45 ;
      RECT 461.835 136.21 462.035 136.94 ;
      RECT 462.38 0.155 463.15 0.445 ;
      RECT 462.38 0.155 462.64 8.665 ;
      RECT 462.89 0.155 463.15 8.665 ;
      RECT 461.87 0.52 462.13 11.315 ;
      RECT 462.245 136.21 462.605 136.94 ;
      RECT 462.815 136.21 463.015 136.94 ;
      RECT 463.4 0.52 463.66 9.955 ;
      RECT 463.47 136.21 463.67 136.94 ;
      RECT 463.88 136.21 464.24 136.94 ;
      RECT 464.535 136.21 464.735 136.94 ;
      RECT 465.03 136.21 465.39 136.94 ;
      RECT 465.44 0.3 465.7 8.7 ;
      RECT 465.6 136.21 465.8 136.94 ;
      RECT 466.255 136.21 466.455 136.94 ;
      RECT 465.95 0.18 466.72 0.88 ;
      RECT 466.665 136.21 467.025 136.94 ;
      RECT 467.235 136.21 467.435 136.94 ;
      RECT 467.89 136.21 468.09 136.94 ;
      RECT 468.145 0.52 468.405 6.28 ;
      RECT 468.3 136.21 468.66 136.94 ;
      RECT 468.955 136.21 469.155 136.94 ;
      RECT 469.52 0.52 469.78 5.57 ;
      RECT 469.45 136.21 469.81 136.94 ;
      RECT 470.02 136.21 470.22 136.94 ;
      RECT 470.03 0.3 470.29 5.235 ;
      RECT 470.54 0.52 470.8 7.78 ;
      RECT 470.675 136.21 470.875 136.94 ;
      RECT 471.085 136.21 471.445 136.94 ;
      RECT 471.39 0.52 471.65 4.315 ;
      RECT 471.655 136.21 471.855 136.94 ;
      RECT 472.31 136.21 472.51 136.94 ;
      RECT 472.565 0.52 472.825 2.82 ;
      RECT 472.72 136.21 473.08 136.94 ;
      RECT 473.375 136.21 473.575 136.94 ;
      RECT 473.87 136.21 474.23 136.94 ;
      RECT 474.805 0.18 475.575 0.88 ;
      RECT 474.805 0.18 475.065 12.9 ;
      RECT 475.315 0.18 475.575 12.9 ;
      RECT 474.095 0.52 474.355 2.82 ;
      RECT 474.44 136.21 474.64 136.94 ;
      RECT 475.825 0.155 476.595 0.445 ;
      RECT 475.825 0.155 476.085 13.21 ;
      RECT 476.335 0.155 476.595 13.21 ;
      RECT 475.095 136.21 475.295 136.94 ;
      RECT 475.505 136.21 475.865 136.94 ;
      RECT 476.075 136.21 476.275 136.94 ;
      RECT 476.73 136.21 476.93 136.94 ;
      RECT 477.14 136.21 477.5 136.94 ;
      RECT 477.795 136.21 477.995 136.94 ;
      RECT 478.29 136.21 478.65 136.94 ;
      RECT 478.53 0.52 478.79 14.115 ;
      RECT 478.86 136.21 479.06 136.94 ;
      RECT 479.04 0.52 479.3 13.45 ;
      RECT 479.515 136.21 479.715 136.94 ;
      RECT 480.06 0.155 480.83 0.445 ;
      RECT 480.06 0.155 480.32 8.665 ;
      RECT 480.57 0.155 480.83 8.665 ;
      RECT 479.55 0.52 479.81 11.315 ;
      RECT 479.925 136.21 480.285 136.94 ;
      RECT 480.495 136.21 480.695 136.94 ;
      RECT 481.08 0.52 481.34 9.955 ;
      RECT 481.15 136.21 481.35 136.94 ;
      RECT 481.56 136.21 481.92 136.94 ;
      RECT 482.215 136.21 482.415 136.94 ;
      RECT 482.71 136.21 483.07 136.94 ;
      RECT 483.12 0.3 483.38 8.7 ;
      RECT 483.28 136.21 483.48 136.94 ;
      RECT 483.935 136.21 484.135 136.94 ;
      RECT 483.63 0.18 484.4 0.88 ;
      RECT 484.345 136.21 484.705 136.94 ;
      RECT 484.915 136.21 485.115 136.94 ;
      RECT 485.57 136.21 485.77 136.94 ;
      RECT 485.825 0.52 486.085 6.28 ;
      RECT 485.98 136.21 486.34 136.94 ;
      RECT 486.635 136.21 486.835 136.94 ;
      RECT 487.2 0.52 487.46 5.57 ;
      RECT 487.13 136.21 487.49 136.94 ;
      RECT 487.7 136.21 487.9 136.94 ;
      RECT 487.71 0.3 487.97 5.235 ;
      RECT 488.22 0.52 488.48 7.78 ;
      RECT 488.355 136.21 488.555 136.94 ;
      RECT 488.765 136.21 489.125 136.94 ;
      RECT 489.07 0.52 489.33 4.315 ;
      RECT 489.335 136.21 489.535 136.94 ;
      RECT 489.99 136.21 490.19 136.94 ;
      RECT 490.245 0.52 490.505 2.82 ;
      RECT 490.4 136.21 490.76 136.94 ;
      RECT 491.055 136.21 491.255 136.94 ;
      RECT 491.55 136.21 491.91 136.94 ;
      RECT 492.485 0.18 493.255 0.88 ;
      RECT 492.485 0.18 492.745 12.9 ;
      RECT 492.995 0.18 493.255 12.9 ;
      RECT 491.775 0.52 492.035 2.82 ;
      RECT 492.12 136.21 492.32 136.94 ;
      RECT 493.505 0.155 494.275 0.445 ;
      RECT 493.505 0.155 493.765 13.21 ;
      RECT 494.015 0.155 494.275 13.21 ;
      RECT 492.775 136.21 492.975 136.94 ;
      RECT 493.185 136.21 493.545 136.94 ;
      RECT 493.755 136.21 493.955 136.94 ;
      RECT 494.41 136.21 494.61 136.94 ;
      RECT 494.82 136.21 495.18 136.94 ;
      RECT 495.475 136.21 495.675 136.94 ;
      RECT 495.97 136.21 496.33 136.94 ;
      RECT 496.21 0.52 496.47 14.115 ;
      RECT 496.54 136.21 496.74 136.94 ;
      RECT 496.72 0.52 496.98 13.45 ;
      RECT 497.195 136.21 497.395 136.94 ;
      RECT 497.74 0.155 498.51 0.445 ;
      RECT 497.74 0.155 498 8.665 ;
      RECT 498.25 0.155 498.51 8.665 ;
      RECT 497.23 0.52 497.49 11.315 ;
      RECT 497.605 136.21 497.965 136.94 ;
      RECT 498.175 136.21 498.375 136.94 ;
      RECT 498.76 0.52 499.02 9.955 ;
      RECT 498.83 136.21 499.03 136.94 ;
      RECT 499.24 136.21 499.6 136.94 ;
      RECT 499.895 136.21 500.095 136.94 ;
      RECT 500.39 136.21 500.75 136.94 ;
      RECT 500.8 0.3 501.06 8.7 ;
      RECT 500.96 136.21 501.16 136.94 ;
      RECT 501.615 136.21 501.815 136.94 ;
      RECT 501.31 0.18 502.08 0.88 ;
      RECT 502.025 136.21 502.385 136.94 ;
      RECT 502.595 136.21 502.795 136.94 ;
      RECT 503.25 136.21 503.45 136.94 ;
      RECT 503.505 0.52 503.765 6.28 ;
      RECT 503.66 136.21 504.02 136.94 ;
      RECT 504.315 136.21 504.515 136.94 ;
      RECT 504.88 0.52 505.14 5.57 ;
      RECT 504.81 136.21 505.17 136.94 ;
      RECT 505.38 136.21 505.58 136.94 ;
      RECT 505.39 0.3 505.65 5.235 ;
      RECT 505.9 0.52 506.16 7.78 ;
      RECT 506.035 136.21 506.235 136.94 ;
      RECT 506.445 136.21 506.805 136.94 ;
      RECT 506.75 0.52 507.01 4.315 ;
      RECT 507.015 136.21 507.215 136.94 ;
      RECT 507.67 136.21 507.87 136.94 ;
      RECT 507.925 0.52 508.185 2.82 ;
      RECT 508.08 136.21 508.44 136.94 ;
      RECT 508.735 136.21 508.935 136.94 ;
      RECT 509.23 136.21 509.59 136.94 ;
      RECT 510.165 0.18 510.935 0.88 ;
      RECT 510.165 0.18 510.425 12.9 ;
      RECT 510.675 0.18 510.935 12.9 ;
      RECT 509.455 0.52 509.715 2.82 ;
      RECT 509.8 136.21 510 136.94 ;
      RECT 511.185 0.155 511.955 0.445 ;
      RECT 511.185 0.155 511.445 13.21 ;
      RECT 511.695 0.155 511.955 13.21 ;
      RECT 510.455 136.21 510.655 136.94 ;
      RECT 510.865 136.21 511.225 136.94 ;
      RECT 511.435 136.21 511.635 136.94 ;
      RECT 512.09 136.21 512.29 136.94 ;
      RECT 512.5 136.21 512.86 136.94 ;
      RECT 513.155 136.21 513.355 136.94 ;
      RECT 513.65 136.21 514.01 136.94 ;
      RECT 513.89 0.52 514.15 14.115 ;
      RECT 514.22 136.21 514.42 136.94 ;
      RECT 514.4 0.52 514.66 13.45 ;
      RECT 514.875 136.21 515.075 136.94 ;
      RECT 515.42 0.155 516.19 0.445 ;
      RECT 515.42 0.155 515.68 8.665 ;
      RECT 515.93 0.155 516.19 8.665 ;
      RECT 514.91 0.52 515.17 11.315 ;
      RECT 515.285 136.21 515.645 136.94 ;
      RECT 515.855 136.21 516.055 136.94 ;
      RECT 516.44 0.52 516.7 9.955 ;
      RECT 516.51 136.21 516.71 136.94 ;
      RECT 516.92 136.21 517.28 136.94 ;
      RECT 517.575 136.21 517.775 136.94 ;
      RECT 518.07 136.21 518.43 136.94 ;
      RECT 518.48 0.3 518.74 8.7 ;
      RECT 518.64 136.21 518.84 136.94 ;
      RECT 519.295 136.21 519.495 136.94 ;
      RECT 518.99 0.18 519.76 0.88 ;
      RECT 519.705 136.21 520.065 136.94 ;
      RECT 520.275 136.21 520.475 136.94 ;
      RECT 520.93 136.21 521.13 136.94 ;
      RECT 521.185 0.52 521.445 6.28 ;
      RECT 521.34 136.21 521.7 136.94 ;
      RECT 521.995 136.21 522.195 136.94 ;
      RECT 522.56 0.52 522.82 5.57 ;
      RECT 522.49 136.21 522.85 136.94 ;
      RECT 523.06 136.21 523.26 136.94 ;
      RECT 523.07 0.3 523.33 5.235 ;
      RECT 523.58 0.52 523.84 7.78 ;
      RECT 523.715 136.21 523.915 136.94 ;
      RECT 524.125 136.21 524.485 136.94 ;
      RECT 524.43 0.52 524.69 4.315 ;
      RECT 524.695 136.21 524.895 136.94 ;
      RECT 525.35 136.21 525.55 136.94 ;
      RECT 525.605 0.52 525.865 2.82 ;
      RECT 525.76 136.21 526.12 136.94 ;
      RECT 526.415 136.21 526.615 136.94 ;
      RECT 526.91 136.21 527.27 136.94 ;
      RECT 527.845 0.18 528.615 0.88 ;
      RECT 527.845 0.18 528.105 12.9 ;
      RECT 528.355 0.18 528.615 12.9 ;
      RECT 527.135 0.52 527.395 2.82 ;
      RECT 527.48 136.21 527.68 136.94 ;
      RECT 528.865 0.155 529.635 0.445 ;
      RECT 528.865 0.155 529.125 13.21 ;
      RECT 529.375 0.155 529.635 13.21 ;
      RECT 528.135 136.21 528.335 136.94 ;
      RECT 528.545 136.21 528.905 136.94 ;
      RECT 529.115 136.21 529.315 136.94 ;
      RECT 529.77 136.21 529.97 136.94 ;
      RECT 530.18 136.21 530.54 136.94 ;
      RECT 530.835 136.21 531.035 136.94 ;
      RECT 531.33 136.21 531.69 136.94 ;
      RECT 531.57 0.52 531.83 14.115 ;
      RECT 531.9 136.21 532.1 136.94 ;
      RECT 532.08 0.52 532.34 13.45 ;
      RECT 532.555 136.21 532.755 136.94 ;
      RECT 533.1 0.155 533.87 0.445 ;
      RECT 533.1 0.155 533.36 8.665 ;
      RECT 533.61 0.155 533.87 8.665 ;
      RECT 532.59 0.52 532.85 11.315 ;
      RECT 532.965 136.21 533.325 136.94 ;
      RECT 533.535 136.21 533.735 136.94 ;
      RECT 534.12 0.52 534.38 9.955 ;
      RECT 534.19 136.21 534.39 136.94 ;
      RECT 534.6 136.21 534.96 136.94 ;
      RECT 535.255 136.21 535.455 136.94 ;
      RECT 535.75 136.21 536.11 136.94 ;
      RECT 536.16 0.3 536.42 8.7 ;
      RECT 536.32 136.21 536.52 136.94 ;
      RECT 536.975 136.21 537.175 136.94 ;
      RECT 536.67 0.18 537.44 0.88 ;
      RECT 537.385 136.21 537.745 136.94 ;
      RECT 537.955 136.21 538.155 136.94 ;
      RECT 538.61 136.21 538.81 136.94 ;
      RECT 538.865 0.52 539.125 6.28 ;
      RECT 539.02 136.21 539.38 136.94 ;
      RECT 539.675 136.21 539.875 136.94 ;
      RECT 540.24 0.52 540.5 5.57 ;
      RECT 540.17 136.21 540.53 136.94 ;
      RECT 540.74 136.21 540.94 136.94 ;
      RECT 540.75 0.3 541.01 5.235 ;
      RECT 541.26 0.52 541.52 7.78 ;
      RECT 541.395 136.21 541.595 136.94 ;
      RECT 541.805 136.21 542.165 136.94 ;
      RECT 542.11 0.52 542.37 4.315 ;
      RECT 542.375 136.21 542.575 136.94 ;
      RECT 543.03 136.21 543.23 136.94 ;
      RECT 543.285 0.52 543.545 2.82 ;
      RECT 543.44 136.21 543.8 136.94 ;
      RECT 544.095 136.21 544.295 136.94 ;
      RECT 544.59 136.21 544.95 136.94 ;
      RECT 545.525 0.18 546.295 0.88 ;
      RECT 545.525 0.18 545.785 12.9 ;
      RECT 546.035 0.18 546.295 12.9 ;
      RECT 544.815 0.52 545.075 2.82 ;
      RECT 545.16 136.21 545.36 136.94 ;
      RECT 546.545 0.155 547.315 0.445 ;
      RECT 546.545 0.155 546.805 13.21 ;
      RECT 547.055 0.155 547.315 13.21 ;
      RECT 545.815 136.21 546.015 136.94 ;
      RECT 546.225 136.21 546.585 136.94 ;
      RECT 546.795 136.21 546.995 136.94 ;
      RECT 547.45 136.21 547.65 136.94 ;
      RECT 547.86 136.21 548.22 136.94 ;
      RECT 548.515 136.21 548.715 136.94 ;
      RECT 549.01 136.21 549.37 136.94 ;
      RECT 549.25 0.52 549.51 14.115 ;
      RECT 549.58 136.21 549.78 136.94 ;
      RECT 549.76 0.52 550.02 13.45 ;
      RECT 550.235 136.21 550.435 136.94 ;
      RECT 550.78 0.155 551.55 0.445 ;
      RECT 550.78 0.155 551.04 8.665 ;
      RECT 551.29 0.155 551.55 8.665 ;
      RECT 550.27 0.52 550.53 11.315 ;
      RECT 550.645 136.21 551.005 136.94 ;
      RECT 551.215 136.21 551.415 136.94 ;
      RECT 551.8 0.52 552.06 9.955 ;
      RECT 551.87 136.21 552.07 136.94 ;
      RECT 552.28 136.21 552.64 136.94 ;
      RECT 552.935 136.21 553.135 136.94 ;
      RECT 553.43 136.21 553.79 136.94 ;
      RECT 553.84 0.3 554.1 8.7 ;
      RECT 554 136.21 554.2 136.94 ;
      RECT 554.655 136.21 554.855 136.94 ;
      RECT 554.35 0.18 555.12 0.88 ;
      RECT 555.065 136.21 555.425 136.94 ;
      RECT 555.635 136.21 555.835 136.94 ;
      RECT 556.29 136.21 556.49 136.94 ;
      RECT 556.545 0.52 556.805 6.28 ;
      RECT 556.7 136.21 557.06 136.94 ;
      RECT 557.355 136.21 557.555 136.94 ;
      RECT 557.92 0.52 558.18 5.57 ;
      RECT 557.85 136.21 558.21 136.94 ;
      RECT 558.42 136.21 558.62 136.94 ;
      RECT 558.43 0.3 558.69 5.235 ;
      RECT 558.94 0.52 559.2 7.78 ;
      RECT 559.075 136.21 559.275 136.94 ;
      RECT 559.485 136.21 559.845 136.94 ;
      RECT 559.79 0.52 560.05 4.315 ;
      RECT 560.055 136.21 560.255 136.94 ;
      RECT 560.71 136.21 560.91 136.94 ;
      RECT 560.965 0.52 561.225 2.82 ;
      RECT 561.12 136.21 561.48 136.94 ;
      RECT 561.775 136.21 561.975 136.94 ;
      RECT 562.27 136.21 562.63 136.94 ;
      RECT 563.205 0.18 563.975 0.88 ;
      RECT 563.205 0.18 563.465 12.9 ;
      RECT 563.715 0.18 563.975 12.9 ;
      RECT 562.495 0.52 562.755 2.82 ;
      RECT 562.84 136.21 563.04 136.94 ;
      RECT 564.225 0.155 564.995 0.445 ;
      RECT 564.225 0.155 564.485 13.21 ;
      RECT 564.735 0.155 564.995 13.21 ;
      RECT 563.495 136.21 563.695 136.94 ;
      RECT 563.905 136.21 564.265 136.94 ;
      RECT 564.475 136.21 564.675 136.94 ;
      RECT 565.13 136.21 565.33 136.94 ;
      RECT 565.54 136.21 565.9 136.94 ;
      RECT 566.195 136.21 566.395 136.94 ;
      RECT 566.69 136.21 567.05 136.94 ;
      RECT 566.93 0.52 567.19 14.115 ;
      RECT 567.26 136.21 567.46 136.94 ;
      RECT 567.44 0.52 567.7 13.45 ;
      RECT 567.915 136.21 568.115 136.94 ;
      RECT 568.46 0.155 569.23 0.445 ;
      RECT 568.46 0.155 568.72 8.665 ;
      RECT 568.97 0.155 569.23 8.665 ;
      RECT 567.95 0.52 568.21 11.315 ;
      RECT 568.325 136.21 568.685 136.94 ;
      RECT 568.895 136.21 569.095 136.94 ;
      RECT 569.48 0.52 569.74 9.955 ;
      RECT 569.55 136.21 569.75 136.94 ;
      RECT 569.96 136.21 570.32 136.94 ;
      RECT 570.615 136.21 570.815 136.94 ;
      RECT 571.11 136.21 571.47 136.94 ;
      RECT 571.52 0.3 571.78 8.7 ;
      RECT 571.68 136.21 571.88 136.94 ;
      RECT 572.335 136.21 572.535 136.94 ;
      RECT 572.03 0.18 572.8 0.88 ;
      RECT 572.745 136.21 573.105 136.94 ;
      RECT 573.315 136.21 573.515 136.94 ;
      RECT 573.97 136.21 574.17 136.94 ;
      RECT 574.225 0.52 574.485 6.28 ;
      RECT 574.38 136.21 574.74 136.94 ;
      RECT 575.035 136.21 575.235 136.94 ;
      RECT 575.6 0.52 575.86 5.57 ;
      RECT 575.53 136.21 575.89 136.94 ;
      RECT 576.1 136.21 576.3 136.94 ;
      RECT 576.11 0.3 576.37 5.235 ;
      RECT 576.62 0.52 576.88 7.78 ;
      RECT 576.755 136.21 576.955 136.94 ;
      RECT 577.165 136.21 577.525 136.94 ;
      RECT 577.47 0.52 577.73 4.315 ;
      RECT 577.735 136.21 577.935 136.94 ;
      RECT 578.39 136.21 578.59 136.94 ;
      RECT 578.645 0.52 578.905 2.82 ;
      RECT 578.8 136.21 579.16 136.94 ;
      RECT 579.455 136.21 579.655 136.94 ;
      RECT 579.95 136.21 580.31 136.94 ;
      RECT 580.885 0.18 581.655 0.88 ;
      RECT 580.885 0.18 581.145 12.9 ;
      RECT 581.395 0.18 581.655 12.9 ;
      RECT 580.175 0.52 580.435 2.82 ;
      RECT 580.52 136.21 580.72 136.94 ;
      RECT 581.905 0.155 582.675 0.445 ;
      RECT 581.905 0.155 582.165 13.21 ;
      RECT 582.415 0.155 582.675 13.21 ;
      RECT 581.175 136.21 581.375 136.94 ;
      RECT 581.585 136.21 581.945 136.94 ;
      RECT 582.155 136.21 582.355 136.94 ;
      RECT 582.81 136.21 583.01 136.94 ;
      RECT 583.22 136.21 583.58 136.94 ;
      RECT 583.875 136.21 584.075 136.94 ;
      RECT 584.37 136.21 584.73 136.94 ;
      RECT 584.61 0.52 584.87 14.115 ;
      RECT 584.94 136.21 585.14 136.94 ;
      RECT 585.12 0.52 585.38 13.45 ;
      RECT 585.595 136.21 585.795 136.94 ;
      RECT 586.14 0.155 586.91 0.445 ;
      RECT 586.14 0.155 586.4 8.665 ;
      RECT 586.65 0.155 586.91 8.665 ;
      RECT 585.63 0.52 585.89 11.315 ;
      RECT 586.005 136.21 586.365 136.94 ;
      RECT 586.575 136.21 586.775 136.94 ;
      RECT 587.16 0.52 587.42 9.955 ;
      RECT 587.23 136.21 587.43 136.94 ;
      RECT 587.64 136.21 588 136.94 ;
      RECT 588.295 136.21 588.495 136.94 ;
      RECT 588.79 136.21 589.15 136.94 ;
      RECT 589.2 0.3 589.46 8.7 ;
      RECT 589.36 136.21 589.56 136.94 ;
      RECT 590.015 136.21 590.215 136.94 ;
      RECT 589.71 0.18 590.48 0.88 ;
      RECT 590.425 136.21 590.785 136.94 ;
      RECT 590.995 136.21 591.195 136.94 ;
      RECT 591.65 136.21 591.85 136.94 ;
      RECT 591.905 0.52 592.165 6.28 ;
      RECT 592.06 136.21 592.42 136.94 ;
      RECT 592.715 136.21 592.915 136.94 ;
      RECT 593.28 0.52 593.54 5.57 ;
      RECT 593.21 136.21 593.57 136.94 ;
      RECT 593.78 136.21 593.98 136.94 ;
      RECT 593.79 0.3 594.05 5.235 ;
      RECT 594.3 0.52 594.56 7.78 ;
      RECT 594.435 136.21 594.635 136.94 ;
      RECT 594.845 136.21 595.205 136.94 ;
      RECT 595.15 0.52 595.41 4.315 ;
      RECT 595.415 136.21 595.615 136.94 ;
      RECT 596.07 136.21 596.27 136.94 ;
      RECT 596.325 0.52 596.585 2.82 ;
      RECT 596.48 136.21 596.84 136.94 ;
      RECT 597.135 136.21 597.335 136.94 ;
      RECT 597.63 136.21 597.99 136.94 ;
      RECT 598.565 0.18 599.335 0.88 ;
      RECT 598.565 0.18 598.825 12.9 ;
      RECT 599.075 0.18 599.335 12.9 ;
      RECT 597.855 0.52 598.115 2.82 ;
      RECT 598.2 136.21 598.4 136.94 ;
      RECT 599.585 0.155 600.355 0.445 ;
      RECT 599.585 0.155 599.845 13.21 ;
      RECT 600.095 0.155 600.355 13.21 ;
      RECT 598.855 136.21 599.055 136.94 ;
      RECT 599.265 136.21 599.625 136.94 ;
      RECT 599.835 136.21 600.035 136.94 ;
      RECT 600.49 136.21 600.69 136.94 ;
      RECT 600.9 136.21 601.26 136.94 ;
      RECT 601.555 136.21 601.755 136.94 ;
      RECT 602.05 136.21 602.41 136.94 ;
      RECT 602.29 0.52 602.55 14.115 ;
      RECT 602.62 136.21 602.82 136.94 ;
      RECT 602.8 0.52 603.06 13.45 ;
      RECT 603.275 136.21 603.475 136.94 ;
      RECT 603.82 0.155 604.59 0.445 ;
      RECT 603.82 0.155 604.08 8.665 ;
      RECT 604.33 0.155 604.59 8.665 ;
      RECT 603.31 0.52 603.57 11.315 ;
      RECT 603.685 136.21 604.045 136.94 ;
      RECT 604.255 136.21 604.455 136.94 ;
      RECT 604.84 0.52 605.1 9.955 ;
      RECT 604.91 136.21 605.11 136.94 ;
      RECT 605.32 136.21 605.68 136.94 ;
      RECT 605.975 136.21 606.175 136.94 ;
      RECT 606.47 136.21 606.83 136.94 ;
      RECT 606.88 0.3 607.14 8.7 ;
      RECT 607.04 136.21 607.24 136.94 ;
      RECT 607.695 136.21 607.895 136.94 ;
      RECT 607.39 0.18 608.16 0.88 ;
      RECT 608.105 136.21 608.465 136.94 ;
      RECT 608.675 136.21 608.875 136.94 ;
      RECT 609.33 136.21 609.53 136.94 ;
      RECT 609.585 0.52 609.845 6.28 ;
      RECT 609.74 136.21 610.1 136.94 ;
      RECT 610.395 136.21 610.595 136.94 ;
      RECT 610.96 0.52 611.22 5.57 ;
      RECT 610.89 136.21 611.25 136.94 ;
      RECT 611.46 136.21 611.66 136.94 ;
      RECT 611.47 0.3 611.73 5.235 ;
      RECT 611.98 0.52 612.24 7.78 ;
      RECT 612.115 136.21 612.315 136.94 ;
      RECT 612.525 136.21 612.885 136.94 ;
      RECT 612.83 0.52 613.09 4.315 ;
      RECT 613.095 136.21 613.295 136.94 ;
      RECT 613.75 136.21 613.95 136.94 ;
      RECT 614.005 0.52 614.265 2.82 ;
      RECT 614.16 136.21 614.52 136.94 ;
      RECT 614.815 136.21 615.015 136.94 ;
      RECT 615.31 136.21 615.67 136.94 ;
      RECT 616.245 0.18 617.015 0.88 ;
      RECT 616.245 0.18 616.505 12.9 ;
      RECT 616.755 0.18 617.015 12.9 ;
      RECT 615.535 0.52 615.795 2.82 ;
      RECT 615.88 136.21 616.08 136.94 ;
      RECT 617.265 0.155 618.035 0.445 ;
      RECT 617.265 0.155 617.525 13.21 ;
      RECT 617.775 0.155 618.035 13.21 ;
      RECT 616.535 136.21 616.735 136.94 ;
      RECT 616.945 136.21 617.305 136.94 ;
      RECT 617.515 136.21 617.715 136.94 ;
      RECT 618.17 136.21 618.37 136.94 ;
      RECT 618.58 136.21 618.94 136.94 ;
      RECT 619.235 136.21 619.435 136.94 ;
      RECT 619.73 136.21 620.09 136.94 ;
      RECT 619.97 0.52 620.23 14.115 ;
      RECT 620.3 136.21 620.5 136.94 ;
      RECT 620.48 0.52 620.74 13.45 ;
      RECT 620.955 136.21 621.155 136.94 ;
      RECT 621.5 0.155 622.27 0.445 ;
      RECT 621.5 0.155 621.76 8.665 ;
      RECT 622.01 0.155 622.27 8.665 ;
      RECT 620.99 0.52 621.25 11.315 ;
      RECT 621.365 136.21 621.725 136.94 ;
      RECT 621.935 136.21 622.135 136.94 ;
      RECT 622.52 0.52 622.78 9.955 ;
      RECT 622.59 136.21 622.79 136.94 ;
      RECT 623 136.21 623.36 136.94 ;
      RECT 623.655 136.21 623.855 136.94 ;
      RECT 624.15 136.21 624.51 136.94 ;
      RECT 624.56 0.3 624.82 8.7 ;
      RECT 624.72 136.21 624.92 136.94 ;
      RECT 625.375 136.21 625.575 136.94 ;
      RECT 625.07 0.18 625.84 0.88 ;
      RECT 625.785 136.21 626.145 136.94 ;
      RECT 626.355 136.21 626.555 136.94 ;
      RECT 627.01 136.21 627.21 136.94 ;
      RECT 627.265 0.52 627.525 6.28 ;
      RECT 627.42 136.21 627.78 136.94 ;
      RECT 628.075 136.21 628.275 136.94 ;
      RECT 628.64 0.52 628.9 5.57 ;
      RECT 628.57 136.21 628.93 136.94 ;
      RECT 629.14 136.21 629.34 136.94 ;
      RECT 629.15 0.3 629.41 5.235 ;
      RECT 629.66 0.52 629.92 7.78 ;
      RECT 629.795 136.21 629.995 136.94 ;
      RECT 630.205 136.21 630.565 136.94 ;
      RECT 630.51 0.52 630.77 4.315 ;
      RECT 630.775 136.21 630.975 136.94 ;
      RECT 631.43 136.21 631.63 136.94 ;
      RECT 631.685 0.52 631.945 2.82 ;
      RECT 631.84 136.21 632.2 136.94 ;
      RECT 632.495 136.21 632.695 136.94 ;
      RECT 632.99 136.21 633.35 136.94 ;
      RECT 633.925 0.18 634.695 0.88 ;
      RECT 633.925 0.18 634.185 12.9 ;
      RECT 634.435 0.18 634.695 12.9 ;
      RECT 633.215 0.52 633.475 2.82 ;
      RECT 633.56 136.21 633.76 136.94 ;
      RECT 634.945 0.155 635.715 0.445 ;
      RECT 634.945 0.155 635.205 13.21 ;
      RECT 635.455 0.155 635.715 13.21 ;
      RECT 634.215 136.21 634.415 136.94 ;
      RECT 634.625 136.21 634.985 136.94 ;
      RECT 635.195 136.21 635.395 136.94 ;
      RECT 635.85 136.21 636.05 136.94 ;
      RECT 636.26 136.21 636.62 136.94 ;
      RECT 636.915 136.21 637.115 136.94 ;
      RECT 637.41 136.21 637.77 136.94 ;
      RECT 637.65 0.52 637.91 14.115 ;
      RECT 637.98 136.21 638.18 136.94 ;
      RECT 638.16 0.52 638.42 13.45 ;
      RECT 638.635 136.21 638.835 136.94 ;
      RECT 639.18 0.155 639.95 0.445 ;
      RECT 639.18 0.155 639.44 8.665 ;
      RECT 639.69 0.155 639.95 8.665 ;
      RECT 638.67 0.52 638.93 11.315 ;
      RECT 639.045 136.21 639.405 136.94 ;
      RECT 639.615 136.21 639.815 136.94 ;
      RECT 640.2 0.52 640.46 9.955 ;
      RECT 640.27 136.21 640.47 136.94 ;
      RECT 640.68 136.21 641.04 136.94 ;
      RECT 641.335 136.21 641.535 136.94 ;
      RECT 641.83 136.21 642.19 136.94 ;
      RECT 642.24 0.3 642.5 8.7 ;
      RECT 642.4 136.21 642.6 136.94 ;
      RECT 643.055 136.21 643.255 136.94 ;
      RECT 642.75 0.18 643.52 0.88 ;
      RECT 643.465 136.21 643.825 136.94 ;
      RECT 644.035 136.21 644.235 136.94 ;
      RECT 644.69 136.21 644.89 136.94 ;
      RECT 644.945 0.52 645.205 6.28 ;
      RECT 645.1 136.21 645.46 136.94 ;
      RECT 645.755 136.21 645.955 136.94 ;
      RECT 646.32 0.52 646.58 5.57 ;
      RECT 646.25 136.21 646.61 136.94 ;
      RECT 646.82 136.21 647.02 136.94 ;
      RECT 646.83 0.3 647.09 5.235 ;
      RECT 647.34 0.52 647.6 7.78 ;
      RECT 647.475 136.21 647.675 136.94 ;
      RECT 647.885 136.21 648.245 136.94 ;
      RECT 648.19 0.52 648.45 4.315 ;
      RECT 648.455 136.21 648.655 136.94 ;
      RECT 649.11 136.21 649.31 136.94 ;
      RECT 649.365 0.52 649.625 2.82 ;
      RECT 649.52 136.21 649.88 136.94 ;
      RECT 650.175 136.21 650.375 136.94 ;
      RECT 650.67 136.21 651.03 136.94 ;
      RECT 651.605 0.18 652.375 0.88 ;
      RECT 651.605 0.18 651.865 12.9 ;
      RECT 652.115 0.18 652.375 12.9 ;
      RECT 650.895 0.52 651.155 2.82 ;
      RECT 651.24 136.21 651.44 136.94 ;
      RECT 652.625 0.155 653.395 0.445 ;
      RECT 652.625 0.155 652.885 13.21 ;
      RECT 653.135 0.155 653.395 13.21 ;
      RECT 651.895 136.21 652.095 136.94 ;
      RECT 652.305 136.21 652.665 136.94 ;
      RECT 652.875 136.21 653.075 136.94 ;
      RECT 653.53 136.21 653.73 136.94 ;
      RECT 653.94 136.21 654.3 136.94 ;
      RECT 654.595 136.21 654.795 136.94 ;
      RECT 655.09 136.21 655.45 136.94 ;
      RECT 655.33 0.52 655.59 14.115 ;
      RECT 655.66 136.21 655.86 136.94 ;
      RECT 655.84 0.52 656.1 13.45 ;
      RECT 656.315 136.21 656.515 136.94 ;
      RECT 656.86 0.155 657.63 0.445 ;
      RECT 656.86 0.155 657.12 8.665 ;
      RECT 657.37 0.155 657.63 8.665 ;
      RECT 656.35 0.52 656.61 11.315 ;
      RECT 656.725 136.21 657.085 136.94 ;
      RECT 657.295 136.21 657.495 136.94 ;
      RECT 657.88 0.52 658.14 9.955 ;
      RECT 657.95 136.21 658.15 136.94 ;
      RECT 658.36 136.21 658.72 136.94 ;
      RECT 659.015 136.21 659.215 136.94 ;
      RECT 659.51 136.21 659.87 136.94 ;
      RECT 659.92 0.3 660.18 8.7 ;
      RECT 660.08 136.21 660.28 136.94 ;
      RECT 660.735 136.21 660.935 136.94 ;
      RECT 660.43 0.18 661.2 0.88 ;
      RECT 661.145 136.21 661.505 136.94 ;
      RECT 661.715 136.21 661.915 136.94 ;
      RECT 662.37 136.21 662.57 136.94 ;
      RECT 662.625 0.52 662.885 6.28 ;
      RECT 662.78 136.21 663.14 136.94 ;
      RECT 663.435 136.21 663.635 136.94 ;
      RECT 664 0.52 664.26 5.57 ;
      RECT 663.93 136.21 664.29 136.94 ;
      RECT 664.5 136.21 664.7 136.94 ;
      RECT 664.51 0.3 664.77 5.235 ;
      RECT 665.02 0.52 665.28 7.78 ;
      RECT 665.155 136.21 665.355 136.94 ;
      RECT 665.565 136.21 665.925 136.94 ;
      RECT 665.87 0.52 666.13 4.315 ;
      RECT 666.135 136.21 666.335 136.94 ;
      RECT 666.79 136.21 666.99 136.94 ;
      RECT 667.045 0.52 667.305 2.82 ;
      RECT 667.2 136.21 667.56 136.94 ;
      RECT 667.855 136.21 668.055 136.94 ;
      RECT 668.35 136.21 668.71 136.94 ;
      RECT 669.285 0.18 670.055 0.88 ;
      RECT 669.285 0.18 669.545 12.9 ;
      RECT 669.795 0.18 670.055 12.9 ;
      RECT 668.575 0.52 668.835 2.82 ;
      RECT 668.92 136.21 669.12 136.94 ;
      RECT 670.305 0.155 671.075 0.445 ;
      RECT 670.305 0.155 670.565 13.21 ;
      RECT 670.815 0.155 671.075 13.21 ;
      RECT 669.575 136.21 669.775 136.94 ;
      RECT 669.985 136.21 670.345 136.94 ;
      RECT 670.555 136.21 670.755 136.94 ;
      RECT 671.21 136.21 671.41 136.94 ;
      RECT 671.62 136.21 671.98 136.94 ;
      RECT 672.275 136.21 672.475 136.94 ;
      RECT 672.77 136.21 673.13 136.94 ;
      RECT 673.01 0.52 673.27 14.115 ;
      RECT 673.34 136.21 673.54 136.94 ;
      RECT 673.52 0.52 673.78 13.45 ;
      RECT 673.995 136.21 674.195 136.94 ;
      RECT 674.54 0.155 675.31 0.445 ;
      RECT 674.54 0.155 674.8 8.665 ;
      RECT 675.05 0.155 675.31 8.665 ;
      RECT 674.03 0.52 674.29 11.315 ;
      RECT 674.405 136.21 674.765 136.94 ;
      RECT 674.975 136.21 675.175 136.94 ;
      RECT 675.56 0.52 675.82 9.955 ;
      RECT 675.63 136.21 675.83 136.94 ;
      RECT 676.04 136.21 676.4 136.94 ;
      RECT 676.695 136.21 676.895 136.94 ;
      RECT 677.19 136.21 677.55 136.94 ;
      RECT 677.6 0.3 677.86 8.7 ;
      RECT 677.76 136.21 677.96 136.94 ;
      RECT 678.415 136.21 678.615 136.94 ;
      RECT 678.11 0.18 678.88 0.88 ;
      RECT 678.825 136.21 679.185 136.94 ;
      RECT 679.395 136.21 679.595 136.94 ;
      RECT 680.05 136.21 680.25 136.94 ;
      RECT 680.305 0.52 680.565 6.28 ;
      RECT 680.46 136.21 680.82 136.94 ;
      RECT 681.115 136.21 681.315 136.94 ;
      RECT 681.68 0.52 681.94 5.57 ;
      RECT 681.61 136.21 681.97 136.94 ;
      RECT 682.18 136.21 682.38 136.94 ;
      RECT 682.19 0.3 682.45 5.235 ;
      RECT 682.7 0.52 682.96 7.78 ;
      RECT 682.835 136.21 683.035 136.94 ;
      RECT 683.245 136.21 683.605 136.94 ;
      RECT 683.55 0.52 683.81 4.315 ;
      RECT 683.815 136.21 684.015 136.94 ;
      RECT 684.47 136.21 684.67 136.94 ;
      RECT 684.725 0.52 684.985 2.82 ;
      RECT 684.88 136.21 685.24 136.94 ;
      RECT 685.535 136.21 685.735 136.94 ;
      RECT 686.03 136.21 686.39 136.94 ;
      RECT 686.965 0.18 687.735 0.88 ;
      RECT 686.965 0.18 687.225 12.9 ;
      RECT 687.475 0.18 687.735 12.9 ;
      RECT 686.255 0.52 686.515 2.82 ;
      RECT 686.6 136.21 686.8 136.94 ;
      RECT 687.985 0.155 688.755 0.445 ;
      RECT 687.985 0.155 688.245 13.21 ;
      RECT 688.495 0.155 688.755 13.21 ;
      RECT 687.255 136.21 687.455 136.94 ;
      RECT 687.665 136.21 688.025 136.94 ;
      RECT 688.235 136.21 688.435 136.94 ;
      RECT 688.89 136.21 689.09 136.94 ;
      RECT 689.3 136.21 689.66 136.94 ;
      RECT 689.955 136.21 690.155 136.94 ;
      RECT 690.45 136.21 690.81 136.94 ;
      RECT 690.69 0.52 690.95 14.115 ;
      RECT 691.02 136.21 691.22 136.94 ;
      RECT 691.2 0.52 691.46 13.45 ;
      RECT 691.675 136.21 691.875 136.94 ;
      RECT 692.22 0.155 692.99 0.445 ;
      RECT 692.22 0.155 692.48 8.665 ;
      RECT 692.73 0.155 692.99 8.665 ;
      RECT 691.71 0.52 691.97 11.315 ;
      RECT 692.085 136.21 692.445 136.94 ;
      RECT 692.655 136.21 692.855 136.94 ;
      RECT 693.24 0.52 693.5 9.955 ;
      RECT 693.31 136.21 693.51 136.94 ;
      RECT 693.72 136.21 694.08 136.94 ;
      RECT 694.375 136.21 694.575 136.94 ;
      RECT 694.87 136.21 695.23 136.94 ;
      RECT 695.28 0.3 695.54 8.7 ;
      RECT 695.44 136.21 695.64 136.94 ;
      RECT 696.095 136.21 696.295 136.94 ;
      RECT 695.79 0.18 696.56 0.88 ;
      RECT 696.505 136.21 696.865 136.94 ;
      RECT 697.075 136.21 697.275 136.94 ;
      RECT 697.73 136.21 697.93 136.94 ;
      RECT 697.985 0.52 698.245 6.28 ;
      RECT 698.14 136.21 698.5 136.94 ;
      RECT 698.795 136.21 698.995 136.94 ;
      RECT 699.36 0.52 699.62 5.57 ;
      RECT 699.29 136.21 699.65 136.94 ;
      RECT 699.86 136.21 700.06 136.94 ;
      RECT 699.87 0.3 700.13 5.235 ;
      RECT 700.38 0.52 700.64 7.78 ;
      RECT 700.515 136.21 700.715 136.94 ;
      RECT 700.925 136.21 701.285 136.94 ;
      RECT 701.495 136.21 701.695 136.94 ;
      RECT 702.32 53.41 702.52 136.94 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 698.505 0 699.1 136.97 ;
      RECT 699.87 0.3 700.13 136.97 ;
      RECT 700.9 0 702.83 136.97 ;
      RECT 0 0.52 702.83 136.97 ;
      RECT 693.76 0 697.725 136.97 ;
      RECT 692.22 0.155 692.99 136.97 ;
      RECT 686.775 0 690.43 136.97 ;
      RECT 685.245 0 685.995 136.97 ;
      RECT 684.07 0 684.465 136.97 ;
      RECT 682.19 0.3 682.45 136.97 ;
      RECT 680.825 0 681.42 136.97 ;
      RECT 676.08 0 680.045 136.97 ;
      RECT 674.54 0.155 675.31 136.97 ;
      RECT 669.095 0 672.75 136.97 ;
      RECT 667.565 0 668.315 136.97 ;
      RECT 666.39 0 666.785 136.97 ;
      RECT 664.51 0.3 664.77 136.97 ;
      RECT 663.145 0 663.74 136.97 ;
      RECT 658.4 0 662.365 136.97 ;
      RECT 656.86 0.155 657.63 136.97 ;
      RECT 651.415 0 655.07 136.97 ;
      RECT 649.885 0 650.635 136.97 ;
      RECT 648.71 0 649.105 136.97 ;
      RECT 646.83 0.3 647.09 136.97 ;
      RECT 645.465 0 646.06 136.97 ;
      RECT 640.72 0 644.685 136.97 ;
      RECT 639.18 0.155 639.95 136.97 ;
      RECT 633.735 0 637.39 136.97 ;
      RECT 632.205 0 632.955 136.97 ;
      RECT 631.03 0 631.425 136.97 ;
      RECT 629.15 0.3 629.41 136.97 ;
      RECT 627.785 0 628.38 136.97 ;
      RECT 623.04 0 627.005 136.97 ;
      RECT 621.5 0.155 622.27 136.97 ;
      RECT 616.055 0 619.71 136.97 ;
      RECT 614.525 0 615.275 136.97 ;
      RECT 613.35 0 613.745 136.97 ;
      RECT 611.47 0.3 611.73 136.97 ;
      RECT 610.105 0 610.7 136.97 ;
      RECT 605.36 0 609.325 136.97 ;
      RECT 603.82 0.155 604.59 136.97 ;
      RECT 598.375 0 602.03 136.97 ;
      RECT 596.845 0 597.595 136.97 ;
      RECT 595.67 0 596.065 136.97 ;
      RECT 593.79 0.3 594.05 136.97 ;
      RECT 592.425 0 593.02 136.97 ;
      RECT 587.68 0 591.645 136.97 ;
      RECT 586.14 0.155 586.91 136.97 ;
      RECT 580.695 0 584.35 136.97 ;
      RECT 579.165 0 579.915 136.97 ;
      RECT 577.99 0 578.385 136.97 ;
      RECT 576.11 0.3 576.37 136.97 ;
      RECT 574.745 0 575.34 136.97 ;
      RECT 570 0 573.965 136.97 ;
      RECT 568.46 0.155 569.23 136.97 ;
      RECT 563.015 0 566.67 136.97 ;
      RECT 561.485 0 562.235 136.97 ;
      RECT 560.31 0 560.705 136.97 ;
      RECT 558.43 0.3 558.69 136.97 ;
      RECT 557.065 0 557.66 136.97 ;
      RECT 552.32 0 556.285 136.97 ;
      RECT 550.78 0.155 551.55 136.97 ;
      RECT 545.335 0 548.99 136.97 ;
      RECT 543.805 0 544.555 136.97 ;
      RECT 542.63 0 543.025 136.97 ;
      RECT 540.75 0.3 541.01 136.97 ;
      RECT 539.385 0 539.98 136.97 ;
      RECT 534.64 0 538.605 136.97 ;
      RECT 533.1 0.155 533.87 136.97 ;
      RECT 527.655 0 531.31 136.97 ;
      RECT 526.125 0 526.875 136.97 ;
      RECT 524.95 0 525.345 136.97 ;
      RECT 523.07 0.3 523.33 136.97 ;
      RECT 521.705 0 522.3 136.97 ;
      RECT 516.96 0 520.925 136.97 ;
      RECT 515.42 0.155 516.19 136.97 ;
      RECT 509.975 0 513.63 136.97 ;
      RECT 508.445 0 509.195 136.97 ;
      RECT 507.27 0 507.665 136.97 ;
      RECT 505.39 0.3 505.65 136.97 ;
      RECT 504.025 0 504.62 136.97 ;
      RECT 499.28 0 503.245 136.97 ;
      RECT 497.74 0.155 498.51 136.97 ;
      RECT 492.295 0 495.95 136.97 ;
      RECT 490.765 0 491.515 136.97 ;
      RECT 489.59 0 489.985 136.97 ;
      RECT 487.71 0.3 487.97 136.97 ;
      RECT 486.345 0 486.94 136.97 ;
      RECT 481.6 0 485.565 136.97 ;
      RECT 480.06 0.155 480.83 136.97 ;
      RECT 474.615 0 478.27 136.97 ;
      RECT 473.085 0 473.835 136.97 ;
      RECT 471.91 0 472.305 136.97 ;
      RECT 470.03 0.3 470.29 136.97 ;
      RECT 468.665 0 469.26 136.97 ;
      RECT 463.92 0 467.885 136.97 ;
      RECT 462.38 0.155 463.15 136.97 ;
      RECT 456.935 0 460.59 136.97 ;
      RECT 455.405 0 456.155 136.97 ;
      RECT 454.23 0 454.625 136.97 ;
      RECT 452.35 0.3 452.61 136.97 ;
      RECT 450.985 0 451.58 136.97 ;
      RECT 446.24 0 450.205 136.97 ;
      RECT 444.7 0.155 445.47 136.97 ;
      RECT 439.255 0 442.91 136.97 ;
      RECT 437.725 0 438.475 136.97 ;
      RECT 436.55 0 436.945 136.97 ;
      RECT 434.67 0.3 434.93 136.97 ;
      RECT 433.305 0 433.9 136.97 ;
      RECT 428.56 0 432.525 136.97 ;
      RECT 427.02 0.155 427.79 136.97 ;
      RECT 421.575 0 425.23 136.97 ;
      RECT 420.045 0 420.795 136.97 ;
      RECT 418.87 0 419.265 136.97 ;
      RECT 387.395 0.18 418.09 136.97 ;
      RECT 387.405 0 418.09 136.97 ;
      RECT 379.745 0.3 386.635 136.97 ;
      RECT 374.135 0.3 375.415 136.97 ;
      RECT 371.585 0.3 372.865 136.97 ;
      RECT 370.055 0.3 370.315 136.97 ;
      RECT 366.995 0.3 367.255 136.97 ;
      RECT 365.465 0.3 365.725 136.97 ;
      RECT 357.305 0.3 364.195 136.97 ;
      RECT 347.815 0 355.015 136.97 ;
      RECT 338.635 0.3 345.525 136.97 ;
      RECT 338.645 0 345.525 136.97 ;
      RECT 337.105 0.3 337.365 136.97 ;
      RECT 335.575 0.3 335.835 136.97 ;
      RECT 332.515 0.3 332.775 136.97 ;
      RECT 329.965 0.3 331.245 136.97 ;
      RECT 327.415 0.3 328.695 136.97 ;
      RECT 316.195 0.3 323.085 136.97 ;
      RECT 316.205 0 323.085 136.97 ;
      RECT 284.74 0.18 315.435 136.97 ;
      RECT 283.565 0 283.96 136.97 ;
      RECT 282.035 0 282.785 136.97 ;
      RECT 277.6 0 281.255 136.97 ;
      RECT 275.04 0.155 275.81 136.97 ;
      RECT 270.305 0 274.27 136.97 ;
      RECT 268.93 0 269.525 136.97 ;
      RECT 267.9 0.3 268.16 136.97 ;
      RECT 265.885 0 266.28 136.97 ;
      RECT 264.355 0 265.105 136.97 ;
      RECT 259.92 0 263.575 136.97 ;
      RECT 257.36 0.155 258.13 136.97 ;
      RECT 252.625 0 256.59 136.97 ;
      RECT 251.25 0 251.845 136.97 ;
      RECT 250.22 0.3 250.48 136.97 ;
      RECT 248.205 0 248.6 136.97 ;
      RECT 246.675 0 247.425 136.97 ;
      RECT 242.24 0 245.895 136.97 ;
      RECT 239.68 0.155 240.45 136.97 ;
      RECT 234.945 0 238.91 136.97 ;
      RECT 233.57 0 234.165 136.97 ;
      RECT 232.54 0.3 232.8 136.97 ;
      RECT 230.525 0 230.92 136.97 ;
      RECT 228.995 0 229.745 136.97 ;
      RECT 224.56 0 228.215 136.97 ;
      RECT 222 0.155 222.77 136.97 ;
      RECT 217.265 0 221.23 136.97 ;
      RECT 215.89 0 216.485 136.97 ;
      RECT 214.86 0.3 215.12 136.97 ;
      RECT 212.845 0 213.24 136.97 ;
      RECT 211.315 0 212.065 136.97 ;
      RECT 206.88 0 210.535 136.97 ;
      RECT 204.32 0.155 205.09 136.97 ;
      RECT 199.585 0 203.55 136.97 ;
      RECT 198.21 0 198.805 136.97 ;
      RECT 197.18 0.3 197.44 136.97 ;
      RECT 195.165 0 195.56 136.97 ;
      RECT 193.635 0 194.385 136.97 ;
      RECT 189.2 0 192.855 136.97 ;
      RECT 186.64 0.155 187.41 136.97 ;
      RECT 181.905 0 185.87 136.97 ;
      RECT 180.53 0 181.125 136.97 ;
      RECT 179.5 0.3 179.76 136.97 ;
      RECT 177.485 0 177.88 136.97 ;
      RECT 175.955 0 176.705 136.97 ;
      RECT 171.52 0 175.175 136.97 ;
      RECT 168.96 0.155 169.73 136.97 ;
      RECT 164.225 0 168.19 136.97 ;
      RECT 162.85 0 163.445 136.97 ;
      RECT 161.82 0.3 162.08 136.97 ;
      RECT 159.805 0 160.2 136.97 ;
      RECT 158.275 0 159.025 136.97 ;
      RECT 153.84 0 157.495 136.97 ;
      RECT 151.28 0.155 152.05 136.97 ;
      RECT 146.545 0 150.51 136.97 ;
      RECT 145.17 0 145.765 136.97 ;
      RECT 144.14 0.3 144.4 136.97 ;
      RECT 142.125 0 142.52 136.97 ;
      RECT 140.595 0 141.345 136.97 ;
      RECT 136.16 0 139.815 136.97 ;
      RECT 133.6 0.155 134.37 136.97 ;
      RECT 128.865 0 132.83 136.97 ;
      RECT 127.49 0 128.085 136.97 ;
      RECT 126.46 0.3 126.72 136.97 ;
      RECT 124.445 0 124.84 136.97 ;
      RECT 122.915 0 123.665 136.97 ;
      RECT 118.48 0 122.135 136.97 ;
      RECT 115.92 0.155 116.69 136.97 ;
      RECT 111.185 0 115.15 136.97 ;
      RECT 109.81 0 110.405 136.97 ;
      RECT 108.78 0.3 109.04 136.97 ;
      RECT 106.765 0 107.16 136.97 ;
      RECT 105.235 0 105.985 136.97 ;
      RECT 100.8 0 104.455 136.97 ;
      RECT 98.24 0.155 99.01 136.97 ;
      RECT 93.505 0 97.47 136.97 ;
      RECT 92.13 0 92.725 136.97 ;
      RECT 91.1 0.3 91.36 136.97 ;
      RECT 89.085 0 89.48 136.97 ;
      RECT 87.555 0 88.305 136.97 ;
      RECT 83.12 0 86.775 136.97 ;
      RECT 80.56 0.155 81.33 136.97 ;
      RECT 75.825 0 79.79 136.97 ;
      RECT 74.45 0 75.045 136.97 ;
      RECT 73.42 0.3 73.68 136.97 ;
      RECT 71.405 0 71.8 136.97 ;
      RECT 69.875 0 70.625 136.97 ;
      RECT 65.44 0 69.095 136.97 ;
      RECT 62.88 0.155 63.65 136.97 ;
      RECT 58.145 0 62.11 136.97 ;
      RECT 56.77 0 57.365 136.97 ;
      RECT 55.74 0.3 56 136.97 ;
      RECT 53.725 0 54.12 136.97 ;
      RECT 52.195 0 52.945 136.97 ;
      RECT 47.76 0 51.415 136.97 ;
      RECT 45.2 0.155 45.97 136.97 ;
      RECT 40.465 0 44.43 136.97 ;
      RECT 39.09 0 39.685 136.97 ;
      RECT 38.06 0.3 38.32 136.97 ;
      RECT 36.045 0 36.44 136.97 ;
      RECT 34.515 0 35.265 136.97 ;
      RECT 30.08 0 33.735 136.97 ;
      RECT 27.52 0.155 28.29 136.97 ;
      RECT 22.785 0 26.75 136.97 ;
      RECT 21.41 0 22.005 136.97 ;
      RECT 20.38 0.3 20.64 136.97 ;
      RECT 18.365 0 18.76 136.97 ;
      RECT 16.835 0 17.585 136.97 ;
      RECT 12.4 0 16.055 136.97 ;
      RECT 9.84 0.155 10.61 136.97 ;
      RECT 5.105 0 9.07 136.97 ;
      RECT 3.73 0 4.325 136.97 ;
      RECT 2.7 0.3 2.96 136.97 ;
      RECT 0 0 1.93 136.97 ;
      RECT 699.88 0 700.12 136.97 ;
      RECT 682.2 0 682.44 136.97 ;
      RECT 664.52 0 664.76 136.97 ;
      RECT 646.84 0 647.08 136.97 ;
      RECT 629.16 0 629.4 136.97 ;
      RECT 611.48 0 611.72 136.97 ;
      RECT 593.8 0 594.04 136.97 ;
      RECT 576.12 0 576.36 136.97 ;
      RECT 558.44 0 558.68 136.97 ;
      RECT 540.76 0 541 136.97 ;
      RECT 523.08 0 523.32 136.97 ;
      RECT 505.4 0 505.64 136.97 ;
      RECT 487.72 0 487.96 136.97 ;
      RECT 470.04 0 470.28 136.97 ;
      RECT 452.36 0 452.6 136.97 ;
      RECT 434.68 0 434.92 136.97 ;
      RECT 379.745 0 386.625 136.97 ;
      RECT 374.145 0 375.405 136.97 ;
      RECT 371.595 0 372.855 136.97 ;
      RECT 370.065 0 370.305 136.97 ;
      RECT 367.005 0 367.245 136.97 ;
      RECT 365.475 0 365.715 136.97 ;
      RECT 357.305 0 364.185 136.97 ;
      RECT 337.115 0 337.355 136.97 ;
      RECT 335.585 0 335.825 136.97 ;
      RECT 332.525 0 332.765 136.97 ;
      RECT 329.975 0 331.235 136.97 ;
      RECT 327.425 0 328.685 136.97 ;
      RECT 267.91 0 268.15 136.97 ;
      RECT 250.23 0 250.47 136.97 ;
      RECT 232.55 0 232.79 136.97 ;
      RECT 214.87 0 215.11 136.97 ;
      RECT 197.19 0 197.43 136.97 ;
      RECT 179.51 0 179.75 136.97 ;
      RECT 161.83 0 162.07 136.97 ;
      RECT 144.15 0 144.39 136.97 ;
      RECT 126.47 0 126.71 136.97 ;
      RECT 108.79 0 109.03 136.97 ;
      RECT 91.11 0 91.35 136.97 ;
      RECT 73.43 0 73.67 136.97 ;
      RECT 55.75 0 55.99 136.97 ;
      RECT 38.07 0 38.31 136.97 ;
      RECT 20.39 0 20.63 136.97 ;
      RECT 2.71 0 2.95 136.97 ;
      RECT 284.74 0 315.425 136.97 ;
      RECT 692.23 0 692.98 136.97 ;
      RECT 674.55 0 675.3 136.97 ;
      RECT 656.87 0 657.62 136.97 ;
      RECT 639.19 0 639.94 136.97 ;
      RECT 621.51 0 622.26 136.97 ;
      RECT 603.83 0 604.58 136.97 ;
      RECT 586.15 0 586.9 136.97 ;
      RECT 568.47 0 569.22 136.97 ;
      RECT 550.79 0 551.54 136.97 ;
      RECT 533.11 0 533.86 136.97 ;
      RECT 515.43 0 516.18 136.97 ;
      RECT 497.75 0 498.5 136.97 ;
      RECT 480.07 0 480.82 136.97 ;
      RECT 462.39 0 463.14 136.97 ;
      RECT 444.71 0 445.46 136.97 ;
      RECT 427.03 0 427.78 136.97 ;
      RECT 275.05 0 275.8 136.97 ;
      RECT 257.37 0 258.12 136.97 ;
      RECT 239.69 0 240.44 136.97 ;
      RECT 222.01 0 222.76 136.97 ;
      RECT 204.33 0 205.08 136.97 ;
      RECT 186.65 0 187.4 136.97 ;
      RECT 168.97 0 169.72 136.97 ;
      RECT 151.29 0 152.04 136.97 ;
      RECT 133.61 0 134.36 136.97 ;
      RECT 115.93 0 116.68 136.97 ;
      RECT 98.25 0 99 136.97 ;
      RECT 80.57 0 81.32 136.97 ;
      RECT 62.89 0 63.64 136.97 ;
      RECT 45.21 0 45.96 136.97 ;
      RECT 27.53 0 28.28 136.97 ;
      RECT 9.85 0 10.6 136.97 ;
    LAYER Metal3 ;
      RECT 0 0 702.83 136.97 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 391.705 0 417.965 136.97 ;
      RECT 386.555 0 388.375 136.97 ;
      RECT 381.405 0 383.225 136.97 ;
      RECT 696.945 0 702.83 136.97 ;
      RECT 688.105 0 692.005 136.97 ;
      RECT 688.105 47.305 702.83 53.15 ;
      RECT 679.265 0 683.165 136.97 ;
      RECT 670.425 0 674.325 136.97 ;
      RECT 670.425 47.305 683.165 53.15 ;
      RECT 661.585 0 665.485 136.97 ;
      RECT 652.745 0 656.645 136.97 ;
      RECT 652.745 47.305 665.485 53.15 ;
      RECT 643.905 0 647.805 136.97 ;
      RECT 635.065 0 638.965 136.97 ;
      RECT 635.065 47.305 647.805 53.15 ;
      RECT 626.225 0 630.125 136.97 ;
      RECT 617.385 0 621.285 136.97 ;
      RECT 617.385 47.305 630.125 53.15 ;
      RECT 608.545 0 612.445 136.97 ;
      RECT 599.705 0 603.605 136.97 ;
      RECT 599.705 47.305 612.445 53.15 ;
      RECT 590.865 0 594.765 136.97 ;
      RECT 582.025 0 585.925 136.97 ;
      RECT 582.025 47.305 594.765 53.15 ;
      RECT 573.185 0 577.085 136.97 ;
      RECT 564.345 0 568.245 136.97 ;
      RECT 564.345 47.305 577.085 53.15 ;
      RECT 555.505 0 559.405 136.97 ;
      RECT 546.665 0 550.565 136.97 ;
      RECT 546.665 47.305 559.405 53.15 ;
      RECT 537.825 0 541.725 136.97 ;
      RECT 528.985 0 532.885 136.97 ;
      RECT 528.985 47.305 541.725 53.15 ;
      RECT 520.145 0 524.045 136.97 ;
      RECT 511.305 0 515.205 136.97 ;
      RECT 511.305 47.305 524.045 53.15 ;
      RECT 502.465 0 506.365 136.97 ;
      RECT 493.625 0 497.525 136.97 ;
      RECT 493.625 47.305 506.365 53.15 ;
      RECT 484.785 0 488.685 136.97 ;
      RECT 475.945 0 479.845 136.97 ;
      RECT 475.945 47.305 488.685 53.15 ;
      RECT 467.105 0 471.005 136.97 ;
      RECT 458.265 0 462.165 136.97 ;
      RECT 458.265 47.305 471.005 53.15 ;
      RECT 449.425 0 453.325 136.97 ;
      RECT 440.585 0 444.485 136.97 ;
      RECT 440.585 47.305 453.325 53.15 ;
      RECT 431.745 0 435.645 136.97 ;
      RECT 422.905 0 426.805 136.97 ;
      RECT 422.905 47.305 435.645 53.15 ;
      RECT 376.255 0 378.075 136.97 ;
      RECT 371.105 0 372.925 136.97 ;
      RECT 365.955 0 367.775 136.97 ;
      RECT 360.805 0 362.625 136.97 ;
      RECT 355.655 0 357.475 136.97 ;
      RECT 350.505 0 352.325 136.97 ;
      RECT 345.355 0 347.175 136.97 ;
      RECT 340.205 0 342.025 136.97 ;
      RECT 335.055 0 336.875 136.97 ;
      RECT 329.905 0 331.725 136.97 ;
      RECT 324.755 0 326.575 136.97 ;
      RECT 319.605 0 321.425 136.97 ;
      RECT 314.455 0 316.275 136.97 ;
      RECT 284.865 0 311.125 136.97 ;
      RECT 276.025 0 279.925 136.97 ;
      RECT 267.185 0 271.085 136.97 ;
      RECT 267.185 47.305 279.925 53.15 ;
      RECT 258.345 0 262.245 136.97 ;
      RECT 249.505 0 253.405 136.97 ;
      RECT 249.505 47.305 262.245 53.15 ;
      RECT 240.665 0 244.565 136.97 ;
      RECT 231.825 0 235.725 136.97 ;
      RECT 231.825 47.305 244.565 53.15 ;
      RECT 222.985 0 226.885 136.97 ;
      RECT 214.145 0 218.045 136.97 ;
      RECT 214.145 47.305 226.885 53.15 ;
      RECT 205.305 0 209.205 136.97 ;
      RECT 196.465 0 200.365 136.97 ;
      RECT 196.465 47.305 209.205 53.15 ;
      RECT 187.625 0 191.525 136.97 ;
      RECT 178.785 0 182.685 136.97 ;
      RECT 178.785 47.305 191.525 53.15 ;
      RECT 169.945 0 173.845 136.97 ;
      RECT 161.105 0 165.005 136.97 ;
      RECT 161.105 47.305 173.845 53.15 ;
      RECT 152.265 0 156.165 136.97 ;
      RECT 143.425 0 147.325 136.97 ;
      RECT 143.425 47.305 156.165 53.15 ;
      RECT 134.585 0 138.485 136.97 ;
      RECT 125.745 0 129.645 136.97 ;
      RECT 125.745 47.305 138.485 53.15 ;
      RECT 116.905 0 120.805 136.97 ;
      RECT 108.065 0 111.965 136.97 ;
      RECT 108.065 47.305 120.805 53.15 ;
      RECT 99.225 0 103.125 136.97 ;
      RECT 90.385 0 94.285 136.97 ;
      RECT 90.385 47.305 103.125 53.15 ;
      RECT 81.545 0 85.445 136.97 ;
      RECT 72.705 0 76.605 136.97 ;
      RECT 72.705 47.305 85.445 53.15 ;
      RECT 63.865 0 67.765 136.97 ;
      RECT 55.025 0 58.925 136.97 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 46.185 0 50.085 136.97 ;
      RECT 37.345 0 41.245 136.97 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 28.505 0 32.405 136.97 ;
      RECT 19.665 0 23.565 136.97 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 10.825 0 14.725 136.97 ;
      RECT 0 0 5.885 136.97 ;
      RECT 0 47.305 14.725 53.15 ;
  END
END RM_IHPSG13_2P_256x32_c2_bm_bist

END LIBRARY
